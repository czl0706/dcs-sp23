//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DgeeoN2sILabbGzXHwVEYWdEaaRWHs7fwdsxwXFEkC2aL1kOUorlxwSsEO+z6uY5
eEDG63VRuS7DW7M1uMk1ank9HymeIGqKLjYqabuuyNTuVuNVUjtY4Av6flr5UK7H
n+RAwj562LoUvDv0UbEwLZm2vRhybM1F7duONmCkQWzDGrSruZjmTw==
//pragma protect end_key_block
//pragma protect digest_block
sV9foRzk2L9YgJMHZDUkfMPup4o=
//pragma protect end_digest_block
//pragma protect data_block
ZDBkLsnYFzja8CKuLbChKL2leTaCbYK9MPeqX6NjQAreOFgeavooljMXtofEfx2l
8Urz2D5RMGGt8mPQdlCEf+9NphPxYeYBE2tvVv//u2WvQ23Dx+BNs4FCmDrqOBiQ
aylzNWAe82YNXj/0Lowdn7KDKpnTiU1Mc8a+vZlONChclzsiTs90nSfPFUAFKhvl
e1KQduM8efFYxIsoauvKmHSwvhFH04+sDrvTUGUaiewWpx9hDwTeJA0drDB9IMmY
CohFc2lvZpDztuPAybnc8qicodYVkpRNU/19mgKDJRfd05LeFj/WGr/1e65PfPJ3
FDTjR2sIihvdHry2TrvGh2qp6n6jPIBYJ+TBCiRovvxgtBTBXuF4bsL3ToBPOmXq
WBkGk5zQ3jDjW1yEvgxthxGWpn0XdVJpyUpbqR8XyC04jcZSc1PCRqSpfw+k4RDM
aDEfeEeU9+8A8z530Pp4ZiLPK0+2U7cqEGEMEUzUJPpq1ozI3q7j/ECCLgy6TwHS
Acy7CMtPECcCSrsX9+z1Cb5LKK+Hhjim5I8p6gXe8OZF4DJcNMh4duXn94CU1npY
ynvMx0TYWp02GvhmxBNKa4RKrXZLj/wApNt/XJH2Z2evlCWJli5t/si11BcKVOMl
RV9gtG5ta7PeKS4h1bNA2mD2nYt0WSNaZ7M6kjJ5O7MvQS/VyKb5XhHajKNDwWdS
8Yh6KXwD0v8PxbnjqANafd7bw/rr2EOrpnOpM72uso3XcE1jAjHPPcvbq9QvGoXh
3KCi1gLJ16myXWxXUpn6ZKRnaIgY/8JqrtsDT9mv0NaOxNL7GsnDqYuYxSkkR48w
Eg2AE/jNcc1zA2fePSqq/g7cLoXxoxTbUFCGV4ydOaE8a4+xL2CwYw63AcrEGvdv
Vzs1iP9rlefO8QFdEhHj3VGh1GjPywaUF6sYR6RHsSOrjYC2IDCycvFQswqIv7PH
kBT1uAuW0T0R8FZoZ5po0eAm67iS3Ke5HnGKLrlo2disZmpUr1IYTlLRXWYyzb9Z
Dsd3fPhfxEzCkiq7eh43SKxN3W2473uhSbII62FJjdycaHMY5T5K9tTzdJXt43km
pqfzXQI3dgdYcK90dJrbhMFxXfdAvTZd4xdVejC8W9hp0li4QxJqoAwQF6hLZrNa
IT1hEcokZh8o64izlUV5SRPpbzA5GW3iXe3uOfpqHzsIk40X7iO2YZhvbBH0OenH
05fc6rGJQe87AunCn9kLZChldedG64Ld5oAffjhtWSyykf8zoe2n86JB6CXxsoea
vjOWX3wO5rZh6PHUdUE6Ee4VrgMqcE3axAfNl91/qv4hWGtSK9TwrSK+gIj9gMOj
emW/8I7BEcsdwIIhvWtLRgBJG2JiHHJzHuAnGRiQwx9efQm+wS7uRWEOSex9SIro
X5Pob/lj4onb3n15KXTjR8+4viYsV7LA+5wYXrTOmCUZj+ka2ojqzA6fNZ1wWlFy
fdxIRI4hzD9j5G5y0s8S2ErlkjFFL39VqyjXyy/MltZB2YP8YieYwPw/qf4dKqj9
EauYo1BJJ4EStcpo5pYRllc4mFzwXR8Tl+fmiNR9A9dMBslE0M+L0IhXwjvziUa3
OT+SKafFpF65QFT1bifx0LBTfI4tbs5mDiIcmRCInaZyt7yS+M6tJTOWk5JRCxUd
o9YXQAdH87fxMWs0qcK5FUBgGPsGUO9Fkybl8TcS7jRIw4VFIzxNC35+Qps8O9Nd
/JjXVq2UJfRq5aVYb5h+1OitwaAPfSZwos1kl52wi04YSDn7qiBaBkdAOQEZifHL
Cil+6pKv9NexLRZV9bwMfpo+K8JUhrfeMKGxWVew8dUZ2AjzYyVAbmW1+g5nSCEJ
1myY/2AzlcwY8zRkSiAW1H7jGCd0p2mzQ/QidAcaxRHp/KNtgmWiXwoZbiS3OEYW
sasaVmnAQQORzCPP+S2nnK/cwh3IDt6AatU0oRaxAZWAIlDz6B3y6r4rD9+MUJlU
vfHIpKFbNEjZgGGIgvg6EKtuBORAEvOm1EiqdBL+LliyjwL3OqrXuiAbT425g1C6
sRQBnBiDpyADuiM3WJlbl1Fu0Ht0vNSNyo6dNq4alid/wcOoQWO0jplkauPGNOzU
YmVSClheLS5fH05shgaldtz8Hrjig65Oe1ujwvCqTVDIEBskiSkn9azt/UI4g+u2
R8Yqei70Fo1Ea/PxB1ObiQKnacXgUWyPrX2GxaDOWUd6erZc4/MPb+StRqBx3hOX
vfkvDYFR05eookfDmshrERhfKOHfAlBd6kBoNA3IDvAy9USY/pui4nRVMi+cONiB
MGE8nxYzTZIpLX7hccifQ9q5cDJ+AUVq9A0/CA/E6gndNyIxZ6JwiMqMwlayb5+/
4+2PgKK6CHIYEqAIh3YnRUVdetcmZ6ii/O2z4owy3fuJHCgf5gWvC3jtLcovapk+
uYGz0nEEDeYdoJm5FWKIa7MeJd13w/FvYvakffXS5/oH0jYl89fO1BOa68HVM1HP
iqj3NYUld1EWsIwMHmtsq55v/dGVF8F/h/CQqosnyXVlr5kYIXwR8E8HvwB5TFKH
DPxLs6KgJGdaAHfKemgFcJ0GF8owQncfR77l/KEftMPMJZbk02p7tbw/UcrJ5yjA
Nk459PgahJ+Kiqyaow+79OByTnfJwfRiOm0n40i3Gl8/ikPh6n9naqLts9uY2Exx
KzCk/jKcUfcsxh+WEtoJzc5DGI772PP1Gy6GGrlICpX/BV8qSCGy3YkdTN5r6y3U
B/YpDmjLRWS6Z9vaf1bjuDo/jRzerkXi9+LxbDvDKfqZjFne4fMHJCOh/fI/lTqk
ur+ik/ptbdlojyqHUsd3QcBRJsu79PZPy9mosA7GaXX2/iteDLJvxH7v3lTcT9hl
vWZ4OUnD+Fglz+55Iz2mxFJ0qFIQiErcVeCGNTXz0p7E3QL5/OwKuE+xyFPB0wSx
bF7MjWRhknSSc4Te3iCELynsCKiSyo4NDMDxHBXWr0S+d/Vnp8hgXkhaDjHP0RYg
chgqI34yWSGd4rCitYkXwiuO+Od72uWJC6U4NtaFSCoO4A5Ly/Z3RkmgJuTPJ++U
joDDfq1v2yHHN6SnmdO+rZrWaW38VDHhMQQVBTRmBo1+e5crFXuZcdBTvz+XfrQu
5wrhaquFs3NRZOHhn/Fs54ORLjL3fNEbG6I5Hl60vR5Biux7WjVSQTsGG8ygEV9g
sBNJi2gW6FWn6cM1Kq46fIxgLuBniM/HmRP9GhWilRIosBuH11lanaVcYCiyphvR
GB36o+WN+SJn/8lNk1D3EDi37MbEQEy+V9f72kx8HCZpqkFuvDXOWV1OUkMh8ajP
Z/ScavgEpcN2oCT0aO4F589hw7jdjAEuAlvE+IxEXszFP4+xEsvd8q26ANzooPvM
j68+GY5/3iCFKbghkgEZ4yR78O6l68ur2OiknjhZxWo/0ZR04RyZuk4SUc7m4ZdN
VtlJg2PFO0DvhkcUyJ3lnSuanVkSxxlOUme4vGJoR7unayPkVfb2vFPVUfq7bO6M
oN5U37q8Encq5Lq6W7R0pel7IPGM4AcEQf7WBdbKNDEW9yNU2E1o46oFlYnV7BOp
ir4BFTW9sdkrulCkxCm2je6pdU7YLUwYW6j9VhGbHhxuvTERChcb527BzFX+5knv
fzZHYNufIUHgR41At250JO8RLXJKx7NG1GZqkN+EXO+Vy+u1p7HXhMNbUFm4hfUa
fNQW73lgW1CjK88uboJtOUiwuY0swen4bufzFL8D9n93ePU2STLeLAwwU+oOUp7u
IznP4ed5MvA6CbBwTvpGkoQGCR6K3oCPzu/5z01+j8NCEJJ74E6ZIuAQ0vEfaeWQ
vJ144QeeVq4bXK+KAIkzGYZ0qhcqsWMuRCa9g8L7YwxgmWxENaPeq8McDZzQlCt6
zegik3/MXb1Heg3IAEMyLjd5DgRwJM0HvJqojUtSEUpCluubc7s0cf2uDkxa0Sw8
hg7oW3LBfN9MadcTBTIbFKxyLCl2jLceDOCjFcfqpi96BQpR99q0ief7s4SUEvbd
TUc+fxVepEdNNhYGY+ceneLUWy8GIZ25dG5ab9m2Jgly3aRIxLIP8dQReWXLpSaC
owhxQrIzB9mA8N2D0Bh1k9Z4FVYI2vZOMKae/7VkHAb+b4H4Xe5S1PTAgQJ7m32i
5D3Fv2cItB7d/J0lXdQF8w0X/gDuq9QgzpnL/D5j68dyoPujwdIrHPWOD1rjgFdm
2Z9vos1eCM/2S3YczynSVtsqGUdyla7LTN/j8ygAOdoLZO0YXw0chgK2Isfj8W5y
4GgV6Gbiwb/qHIWSsJ0xs8tzIZo/wOpwKgOsfuhQk3Sm8rHUjFSmWPCJu4XhpEyc
NdtImA9j8+9QNyavCx7cSwDpave14TNyXtZYU3ptOPCi73tTPDc1+GdOOnXS6l6f
3WhnwZgINaiXu2zz7Lh+fJaCwuGra07E7Msxw+4JuId0/dJpXUnAwdTL2R227aLE
89YfMQg91+7n8Nj/Lf9KJHZ3hIrdtrF/qNwfAjC4xB1ct3t5zChKFqvu7lzuMPjl
nHW4N696eO7t6Du4coMt8QOg4O1eDfdsjqzbVFDDknAU8E0i//Q7w5JVE4AFWSwt
VrZF/zcpvpP+EwKCBTFcKhsBGEplfjOtlxulHJsUK2wEZbwHmj2ATkLJFyZo5/yf
hgDVjz9lhuPWdwMYsjA1W3UwuUM2T5ueuBM/1iJJfmXKshM3rp8t5ooLqTc94LGm
ri8RGdAutfaGSt/t4Jve05WYRfOgY0cQcaLNJFDeHZRm2so/dSfNw+ZutRtN1Bac
VeaQIj1A1Dzwy5McWwu6n/2Q0Fx278p2BemFDZBTfbaISpL8iSL5sN9aYGjwwcks
N7W+Ag34IVL+nbbbTcLGNjlCrfSjxWweFe55z4FL7Bj9a50nF7w+3HtmpLvm9l+2
znFeHI2DB19rhgTlCEaVnwL1TDlJnGbc+HMNbiaWP51awtclD+Ize23Sub2Z2SCs
A9nJFkRJGISSQSPcNqh1HF9QTlK6kOljyDdlDN7M+op5kGPtst6fq896qhHb0LHi
q/TEI09wIdDoiHkliftVen6W9TXhPyeTK8TMqm3aPg5sUKHhe0B6Or+iA9r6bNsJ
sMEGgcacZaJ4j/Nlwxcy/chpKnFVq2bsIfxnkobiR1iMoMGl6xTi77+Oqws+Z9pH
8ci9fLP0ePo683ms6ZItfgaWPckB0n4IAnIym4wswrUjf9tv1sicDyaNA8qLqQ+4
MEXGY6mxF3GHLb9ySS1vjIhYgVRvAL+WnII68ajAvJIFl/TnA6sDQg8GFOhY+kMr
4yyfZSoIcHBCANdPjZnE22p6OTrJQ21eneN/D8kGDzyxc+v8+/qZkELbVo/FE/fp
wkLDsIUVuA6abpzcAmj0g73W85uXlYWtpFLldcVleLDxu5YxEpi3KAL4B6BXEg5A
RdJZ6fq9Ck9rTlLtuoNyCqDQLDM6Dv3KIqYLipR78UTsRXODTiUvO39BcgugBLzf
5t/PJQDJH+eiYWuTDw8eOWMG2hW/+brDZHX6gHV7nN3c8NTC2mUbknKVh2SMFx6+
i4w7tgaOVJthnL7F9VYuBD0LuvUwGKRBmxYtDMKJFXmXRlm4PSf2knCbiGUmXcSq
ykD/OG2PHvwQIkN4wICtZso6TPDnFftcnTPSscHTkxphhlqaJVDZKbpzHrPuCHAR
VmwzwZdV8CMyNACVYpwxBo/RB0OJdTGPuQtOn14mmdepduSL7/W6VkLRhD8OGoj+
cK8DsQuZVwwHjdqgPBYTFn5FjdJeuN9XOrykPd27yb/oWjF3r+ZNquvvbZpf39ai
zg5Og+Gcvg1bGw57BGENU78n8hHbAAoKI182wfj0zYyFZnx16aNjXizLiU4qgBOk
WLPRYjy1rtI30Gdftp9HxLmwYT2odAkIHE3iC4lF3xn+F3n5tFwJsbWWB4M183iB
FO/TYneYHpAs1Ki4mhC4HiOd4Eit40ZYcsTj8V6i7gw9+RvEemvT41w18+NNlEUU
8uPD7xUNbmvjr6WvsHZ7XCQ3TrCQjjflShTKZ4Fld/AnT6u660rf4IYHTOU4lSGG
CUG/8SG/MlRAYI77gpEPsuvNQqd2YZXQnKvcOcsHFWRuVWh9eUZWYnBuYUMKW4xb
XQ53YR2Oq/DD2NDJu2fln0nkkxR2NqoXCgoDsA98eQYzR/O8fxiC2vLX+VdH/rcr
oaIPg6YSmQKGeXfC3Pw7dx+z1vdHms2CiUb4xrmlsmdLpOYQQEmPhw4IN4iKxCls
+uVfAaoe5sRJZH54ZBbYP1K3Ff/ux8ih3t5GXrpKFkNMgjPMm5bQVeRY1hBC2asm
1b5Ymccm2DfV08EFxMIf6aa8EOI1/IZAbd4VqJGSbMacbQyKn0DOvcspnFPyH21e
Iw8gmRNhkvdcX7/a7VAHNLQ5wOiMmo4Fmi1SjAk2Q1Gm6DZ165s4KYK/1OFi5mp3
s4OMjJ90ai6LdnJZFw+k2RJvh+hTsdOLi77I6dE1YoniHoUUEyA2okNV2cIgnrrx
T16szsvZNTYinafv7IyCAOKTNSPLMXx5DhvVrKhlNlGW4TmxbHFQh9GsAKXjaTSQ
xspLUxwZ5DmUUAFZojKcHoZCScBnHPiIB4xjT9tl7lt8WsXtLIiQ47Vo8xiN5WKd
sP4InsMuvbLzIF4V2WKK0Ut9L7TUIy+noW92xWSYZhKJvPScTYvFvaoSazlJ8qo9
lL+XI/TaA/+N6Qcbh7QX1wSHAS+XkXjrddFeC1l2HRDF9E2ODyGW697MGXB7NAns
1uv8PEhsbWYtjZECG/jXPA/Ha+jvjjP/zZxXkppLts9ObnzgWIUMktBcjBC9PY1O
LNdAKkKa5JAeajMw7p27MB8wl54a5/7TH/3CHu0rz29VJGW2F9O+3EdIOWIDb2Ea
uWG58ofyYzsLCp2209Fh8FtzBtZNGXy/b7MGbbMT9xqiFDogJNqjZBq4UXUW87Is
opwxxvfE8Er2UZJnhkMmjVy1LGcGa9ew7wXGwULNpNZq/nI3pgtPHW0eIQaGdcmX
i8nfeTEXyuEu7GZRPZikwURxtov0qoVLq3m29frIXygWrz5XPe6OKEvgKYBj4bpd
BGJN3OsKVtV70CEe52lytgKzooBgwh78J2E75omVRxHQRLbMGCGACTD9O8d5fhQI
+L8s7D3KqSXPwDWsQUvOfxidOv6rgy6dyAocQIcubxlucg1VFt4txKSJ2gicmmEJ
EPJDl1J30Y3jTlxe7EemG1ZLZNHT9uPKTiFJZnzO/Ij0GjCZfHHnBr8y80Ne9ICc
RxDTGA2MrYJ8mQhsu5J7GsgMF9s9VtL+Fn7QfdwYi5u3xgHWuvQe0yzOzEBvwx1d
TunVqfb/SfqJzwBUlki+JrEVE+zLu7+m2ylxqrVvcaL1dvD0mvbWreq8+vFCrADv
6nTxSO9l9WFTaX0bzu3IJhpSrc1ejfcT6MwPjbDMdWQbdNRTnhCa7jkrlQHvJEa/
G/S4cSmFKVpmPrZqx2yEi2IKgojf+A1p3y3byV9SGYhZaRyTnXrszrTKG6EreJkp
vtT1xHcOyPp9PSoSgqvTYgzRGlW5ImFQgf4LyZ8kdvTFWjT+lvTNWG9upuOumx43
O6KsZ9Rbv7lw7871dJqLKqpq2TavwMaRKHqCqMVvlUxqK8Xy1cA1XvMVaMlUmZgL
BK2Qj3FsJnEUjLL2CMUbWxLlMmTxYW5UxTXYx9b6TPRFmivbvLk4+6Rh2FV3w8NY
xvDbQwu1wxjnIKmc/7r8hGmN4vWbOB/xVv0FkS7IvGVzaJCgTKQmMGlI83JGImEk
U56avqDs15uFRnfs/qOuMYF+38/VIbfxHOlScNQZGmON4/QXWZirC27eIOJ8dEhx
xquGEDV8s7DfzGjn1Mc7JoqrELQHaE2gKo0DD7OX1TEm40Er9xkJgTAPhyiAXpaV
bqOTe9p7iBuyFsGP9A26WJmhtdhKg4sF2DuslLxiLknaNGEId830MPzoOUR4PmLP
RCuOa5RtAGYgRiJDZyA+TwKgR55eM3Wcu2J5A+QUTvdpXLGtw66T0kfdiMMOc2br
+wV+/kbeZrWjv7aG+pr3d0esV4kByv7Y9G5HuQZQHUKRS7UE1ojfhScjjin+aZFt
k4LEmUFx8Gr2GJV5IQqfEHLMSJUyLNYA9Q6As1wriJXCB/nfFfCCrJloAbmIHFZg
mnMOj8UFhEGl+n+I7EXI6dK/W4NNlgkpscpOyjULnXV2VJRaCT9qHVpLNQg8wfwE
3m2E5DCXFGL3VZErqKvr6EOMS0CPUc4nwlt1brBWMgybJaAo8QdPQgwY5wGpcIDx
uWD4e0Zvahg2CUQnaBtoIlzfhy3Lf9Ktu2ENAePAfTQTafqVF+TSaiII1TrNuId7
5BJJ0iED526FZ15NtwHPmFKb/MRfHKL4VyCH9iRYyFkrET0/ycrF605fo18m9tQb
ZknQrV+AkqASFjXywXMSiKLRvSO5NayM3KSTON4yhhckDxfkILzIBihYUTLQ1K7p
zY7uiagvj0BSYpdKbXcdiNw1CfJ5dB4KRc/jOmPSo2g3pGpYmTMUXek/dkVJS6at
gKsHIpAmSS3DiLoK63imTcAL9DJu20ICQZ6j+Rj/Yc24ojE4E1FIOLVkmA3hHkWQ
IUN5nzbHxYFpoDSTYi+kuJ0oIsRJZDQoi2izGUqsBGeUp5fl3QceJKQV+p/Y/ZEF
qCJCG0glxyax/VAfU5sJuVAUMVcdBsXT00W2wqI3F8oKWUWzOHbEj+iwrT19rf+9
5b9H1AW5c28jDwh5aVhPSuqPJUZtIwFe2ZMUw+S9IiD+t+FkGDSFde9w5uNSfRgh
wSdhzxNS6TYxRoXNARLYh8R1efDH9ro4vXnK8U3KPMI/4PwDoeKPb+jsTPBclNRA
xyv6zi53jU+nLxOIYauTnbX84H4QKmb/6HEtPPWhxpPk5G0zCSN1Sy8IURG5TCam
zxp7oGnzkMz8ftzaTPpLFc80pm0t33jvhZVQ6pE600sDAZYs4ehiUiwWTal36iLf
Y7FCEykAJUm0xaJwlQcDrApj5RXPq6c8J7xBJYFxT/HqX27TycA6RqLL8FxKaHKI
k6pW2jDnqGjriYh6/5ZSkPTlbBQjbv9UtfJCB7ab/kFB9gqEcBwAjJp8Yy09PmLH
XcvGYCnlXeZ2nJ1l5Rk9c35Fe4qk6mNnHJxUFEnJ9r5+6hffFUmLs1WpOJmZKnzR
FsRcvJmrCaj5G4RMQXGkWBgKX4m4YKYwKNFsak7nJtCOxMbqo/1cXUx18meToTBC
7PIJ7vbUY2BDQg7SeZE147w2MMosAwP7MmfwgHkykPzF5QpIitQ3XKOA7UyHm/Kw
PkBENNWOMqULiv/7ezbTI7Wj6ctzOt2kDUvr0bODScnmWKdZH4VybWZzkommPIBN
SBuinDKwuoogWrDsImogweBQY9L2+oFZ1PcTppZZ2N9DF4VCDrn7pJN5a6Wpjk2l
b2K4t55029+X7r7NeISPVbvFC3lRwj32BSAAok8G0wodOHAjpn+8FQTdzcq4bvNF
TkyH+5VKwLv+3/VVGFkTG2/YrA+cV5yDvq9KbwXBo3D4NCAwHnI8K/w6auoy7iDg
LGAFNVdQa5L68qCrKeAgSzMIQ7Me7jglMI8y9PkRAtN3J7LDWDTzrQstV1awCoww
Bo1uKsvrFCSNc19W+ati6ugDmxM/LkrxHddbBTIr4q8cd4cIxgbym0JTpR5FMw1W
Tep7xuL+nMMxDvf5/jju3hTloh2D8VxU/VkOcHY8OAWInS0XSZVeU7Xk1qqZmBJb
CDJdvO/OGdamvnETiLw4bhJ0BGPkiGQSic4336KIBqym1G9+Thb508MKVUjKHU3Z
eQSk6eLvFc5VxB49r1Z903lLLn3V28SZV085q61ub3oD2aqVZh8GBS3ACGkRpzKZ
ejsIEA3/6QT0VoDjwA9Gk+oOXITtgu8MMZK/el1peKl5rst6d0Mjb1PxxFdxqjk7
7DIDmpnhbRu1aIUpmYdNCdYTYCBZvM5GShBoXAS+edt1mIBiB/ON4lCEYIW9KcTa
N7cva0bmtsGKA11Wy//2xa0P0HfMyLHUl7atEi8Nla84Isa8+hD5YeW59X3Fvw9q
7K3LZsID7vApXeNZD99Dcbh5g7fkcr0nUPTdgMHZlfxBIoW6dgDY4nCJVUF5NCJr
DsCm30hBp18vYP6r0/+MtO7ibL+ZIHr2ehIrEtaz1saH0ZFPBimbWQHmdt2+PL55
VeZCVD9JTQcO+KusRxUuqJWzcgTXZbNaJZmDB8LrrAKghPKeweN8V2vqruufQcZN
PMRfsyIfUy2YRFxcavim0Qebkc70+nS7vUvjBaDCeQfMfwv7wPuURBmIdBGVMnTR
kPp71qeqrvov7SMMHCac9KQqJj19P7lgs/406qcLRiL01gFpO1NMehnlnBoxSXiC
3DOTM3mnFKIkp44KPkHioy0x9FajFCBsFtgKjHWqR2bP3n+w5LPrKu949n597wHu
e515uip383GnFwsBQXWuNbYQdYAzkrR3HRrVlBGHjN6g5QLoxRPwsRnpdADP4l97
9eVpt+nsOuFPdw4DcWGk3KxJbTD5/ENJ926Fnb/bpKdLXGUXAyYU04o2Yy6AbGgo
KCTeZFSzp5Vbg4c0y24Hcp1CscFTSD9IVyfyJWCFsv8xbaiQyjR8FtU7HVW6dWhg
nS1eGDXvdkLgr9ECyBEJa9QuudDQoAaVtyfFee9s3Lwr5M6H/PV3YvI4Us/dgUxq
KTR4fUyCMc0lXUasJioeMUL1UjRTLhK7Mj8OoTyVmaI2ClNrpnv8oYNj2lRkAc7f
JYBZrWMWEAkva2lJUFFPAToVi0TjFIVSBqfN9H2ZptqojUHz7/JptbEiaTBLF54O
NkUvh2Jv+mS8uMt1nANQHkqqVEqm5w2z/OcSySjWZ8zUxsUeiaEL7WmOApIsGRLk
CptblwWoyHO69QVZCxl3GzX+LpcuESQrWiRTerKShExxmFZZX/AeiK3MqpqvMXgz
F4ryEKVTGcDeki/mMmaCb64EYnIeYRxUBtxN6NCFTrrtov3IUcXf3ur8WMXrzepM
ARTnUKXhHEY0fkocwJ7ECe40GmmnPVuhDQmJRc8WbcdjGfKxjOWxmED9KE7BwjZH
ecLETXvaiDzFhWpiCthIVrSZHDXN87/mV+VkClw6BX45DpmNVDuWC5XV2qD7sMr+
Pnqf5RWyGRVmFE7hmj7zMu+GuFryjVpm1pALJOBLyyGbfz4Tl6rFA/tfqAdqotRI
8pGDQHCUWgE/bpShdoU/tnbHhS6s0amB/dlTwDra9jsdfLOuNXcZapD72E4NqvmW
08vF3CJfAfC60IAjkB6065pQ76LAisato+v4EvM1dNTfmBinG2mt8rnoOg4yI1Gs
lJctoEerMouJkssD1t1p1q+q6uLmNuv3scYIZEqaMeAK1kq53o7nqDvBmhcmFD5i
83IPok49nq2eXmKPyT+Br0xR+tKtp2b1rnjJdLy/4xZ6eDV7BvbxFt+znafY7p1I
cOviwHkM/Ts+fLlCVM881qongO4FxvImt2/iMNWB5B7UKKE2cKWvaWPxAS3MouJ3
8vUFdOoaTKohwUqIcFjS7kAjotoe/MTVgozzL91iYdHd/laLbU8VPNx6q16GiJqd
FHSL8uBMxWJYi1Ao4QWUcFRZj7bWXtVPI1GlugOyf/hxGpZAICh/0yyNfUPsesJm
r0DnxmXGSmhKepXReWLt97g+s+lpIzgZBxZJLJbfZJmW62t59XhY8Ws1RNff8Ei9
cjWfOawFq8i9tmJtB5usctp1OSWkkqkDIaBW9hfvsmjnqYsT174+cv+hup5yDphS
KBtszNeVet2C+KGuIw+5Dh9iX1Z7ZLI9FXUGQe33mnoVSMZO9/N2TbdHAJZwBunI
auoGaW3gW86oEPKChQIXZlvkqNW3UaVNIPMF6lwOuA9ZDHIA75W7/Kae7qxgCDMm
StL2DNrmLshmLXo20hURWutXIAYxRT0Ro89sgG9mOCZPC1nv3m4db04DGMpuhKrE
P0ncxeQOxMLE4WfbP6F2ijyUOqxV3y6UCVI2jVUlijT6yrdYfcj+K6mqApJqFyFp
OF5+jBYK18bsUS1fR/pEEcFJESj/ZY0T9bi8iBdsysX7tpTpFASqf+aDtVhA9eji
QJqd+LRgKuE6BwIuDvZjOexnF9LGdTSQSxJJg3VrRdYmhSrrnqKXfoQ6oMpjlZom
V5umEa3dRLUovg/ewciFEmtPD1soH1bASF9S8ow7W73bK/+9X8fNozczJaFUUGS7
5b7x5BssWnm/xCRvt27DW1jqAsdqT3OMuAkz1TpQMKlizi2np4RzEYNKBMxhufR5
u0QOqIczXi2eoXBYXBKYUqC+rp9tRPj9zc2fmFQWXbVOphyBkE8Xme5u0za5Qo1r
5WvltRkYNFMO2A41yU5vzieObMqFGxS0kB1R5rHDtuEExS1GGSvn5qu8bwO68f58
LgPWP8TtBQd6mUXE0ToV3zpm3B+4UdYvz/fEvUXTvxfgyIcvN3JdCFd+LncmV3XJ
NivY7V6LB2yPk5AalBFGjdUPdAdcQZFJWqqJZ0jM1vLIOidZjWNTYgO0C9vZw2F7
Xe8LclB3M9E0Zi2iAT6N04rPP3lYoVo39WNeTv6SxGih8WcSEDTKI4t3wf/GStiu
dKcsQKRCkCkiOCD7xVFdxsInSShgySFaSaE51Pj/2YWwK7dYbmAUlWudSYLPofSK
ntg6mCxxHnBtH9/lwyGnbsXtGBOpWbnnAmfGUQYJPGjDK9mvzZUHH+4tH00Vu1+u
ZTTRFRihMChNtLmOnuq9zWx7OLS4Yz09xrQ1XG4BjfLorj4p26RgAF+1qZ9mbOAy
P8QHR7unvSoFI5rCCPUQIRdwWyDrz0/5UOznprXrZOrA2FEj1ARRlBuv2TS18NSM
tV4A92FiDneT47nKHJkJQM/qCCyoVzpT2/d5oJjKUeBH2IhIN0iMS3AGZLfvGJeK
SdrE4FMQrQZ+Q5H58ZbWzPLRGcVVtNQKExsmCk8zE0XNqK1Srd+b6E25hKGEyXFZ
5IiLo2p+JOBoK+EZEhn1gIhRWzNNfgDvvT0hajnA7g/JKcbUsMZLTo+RfgCKycei
2xBx/WO9HUtNk22oS4zWa57wuizubWhDf8Sf5Eww7azFbHsbfUdV006ifxPOLdug
sRlRG++2bTxlgKbFrcPNlDRGo47uv6hrGCNb/xIS7wbsn7UHeb6rMsDOq32e9dX7
HPHw+V8Zb/klOARnu0hG/rlmqkGACVPhPtnhuwyyqs29MmszduQfenyVOCYVr2Ig
V4UHaGP92aWiFiMzr85hvMocpJSJjz2FLLDF3n+v28vmZ+hf7s0Uo9F7fhgLHoJ3
wGzpgs8HNPwB6jzlAtaBSfsxCEfk6pMo+s8YZZVkOgGsybZOSu5OaGDdI2ScDxS4
ebKZRoXTCiefUrO6bg7meMOSksxIsDlSbPpWGtdL3Ro3rbYoLj80J05R4epDJHfh
veOR00eLRIv8kDjdAbSFOvEuX0fky+N+jfXcvgGPCSGo1Zpz3ajd20O5Od74Wb6W
iHQjDBSJIzVQY18N3mR0CSQe8w0InAUR4wc3iR7Pu+SDtI21k5pcKUmjOr8e78if
kY99WjmuVPzrl8uTTigRXcsjmZnRWSM4OfthsUwMiFTQ9R4pREZSbClcjMRLHFrP
+APKsThmtRzdylfJ6dUB4O/u0YJZ+kW0SEKMYvkH8B7oacrbK3b/n45gu8PTsrIl
YzMWRzgNoYX8ofHx3gSJJxT7ht2OcG1HuzXL73uIy93kC2OK18l758v66AK/2z/T
pBsB7N+Dwey4TLZbkuD7hAdXyLMfCK3EAlSDE83+bRBdHhJxOrqdbsB+t5OOW2Ur
Rr7DizKz2tCdlkU1oPUK1vxabClMnhVCN+PcOhyIFmkfbsVjgqROo33HHOYcpqQ/
7uPF0/v5zSNaqZ3WNIDO3VjryfOWeD70/7JPKcNlmDLuhjJiaj/7F8ghwytx1Owh
SpXfrLNXKt43vpwSmN4pfHDvB7IB7u3WK4SktjQGz4vFv2PL/0kcYJOj8PTPdQO7
QsXoNdxpSlhQRdYXcua++iV0ipMG3fb0NdM1qv7ERxcz3nqNYhZSDSfn3qX6xeI/
S2Ha/DfF3l/jfqufeMnr+/gLYTa33FPEMYtaox25C3jgLe8x6ykhjebVE5EES4y7
Z/dbE97guyElAHFSqKHU9jBX97LOYzS479dkY2LiPSjdCfM8Lt7guq/hz/lZnwP6
EOw92AXDIqmfrghCwIqDEdyyf+awYLl3SFkLzzjZQVy4/mmouDfCRg21vYY2OX4I
AfXIkpzoFNu5+j8v2jxrO8HZs+dVlE9N1u7VM0pe1kpXGPCSQodnBo7v6ISz9/VH
M5BpdyxMnNoZ0ixmP0zS55diITQOUuPjPoFrz4HEv9x0OodfBKNf3Ru2/6ZNLhix
5fu278zbbXpBrhcyagfL5TElZrkJnTYbf4eKArOpFKCiEfdNOWPeT/NfRfZkUqlW
LJviOa339HW7aPtDyONvKmEwnM1K673qfMJWW1oeW2u1oQ8vM+v7gsQ+PWbUZBEt
Ef7GIaYGZaM/da1gvYiMqS66AHOdY1l0QtDpOitBFVpo0EDslTRCNYjp10FRCv98
hWLV/NazBlD6rMFNTegTNP9Rc3Eh/6ymqJgveg9jCADEoEPktqlfxgqObdOcrvKJ
B7EN+t0rTAaGe3ZeJeXqBwoENqaZ9sIS+1v9xV/9JqkMTrPbvxsyKnfr60LwBAqu
S92w6/WOYSywuozn8XgMlFsuUTQti1BrOkt8IV3fF6P9eSPorYGnAt1Mp7VSa/S+
LdTbvhXUnCODgPgJqXNfUoY0Lc1TwQoF3krIvbzThX73LmCAbs8TflwXdsAZRRYR
zyg5aHqpX2vsjWGB+cxT2ZS3N9Wo9HCohtvVD3DM8MeQjlkIYU1pp6C96RCgjkbQ
hs50OzErIy/nVeF0uq4D6eoy9JLSo03Nl9nrNVgj4hra92s/se6fA25BedUEEX0s
MWP0cMyM76eIrjk6JCZkDi95usowqo4JKFDMMQpKUxcaWBqqYC7MipE2JtigkmWS
tNh4mcYUUmoGUOrRi+qMZGMtpQPP0xsnXBp7ZV7WujbzQC0Bl+UIItJBs2KCJfg7
01PmKbQqPQK1L9X/uJm/NSnE5abFxiVbqufDg+RTaA7SvVFjFhC5lEMXr8rT05Ab
4khYd9YpDj12LyQxnS0fgr9PW2KIey3He8H9c7EggrqLlaY8T6TbLWf8Kg8O0fhB
jj76idlMTtQiGFUq0mWsq5zM/NIWkHW0ZS5nE7sb0YyCFXkKKNYX/uTVRJ/B13oL
p9m6Rxl9R6PH6zktq4NinezIbNR451FTYoqtLys6NDNplDQDKby6/JGhRKLMjmLB
fgJQXrDmLZCMbEEVqXy2bL2jTuZv+GOW8JYUtSt5fRiADFwn/KB0MXOrOpnwa7u+
Mmnm6YLnip0Wuh/LmqPJKPPRbU5VW+VBDFALgZDipT8Dp8JZfGBSnA4RoTeoBOYP
iNtKmNdCSCDYg9KvZ3v6FLzemygtDqOgSg0bAkw3fzJw7JfcG4MPjICUMhoRp1y7
VzCTg4uIYxbrUkBlSVJjHNYsponfnPcmQIgBYtogbfjOctVaos8o9Cvvl3fzFg/j
T81yLKOMoG7HzTFZsdmE21TfgS/EXwsbQmqVWmFk1Cvq4FDMdwCRNyoEPbTD9FPU
9fvSFB+vuZsEXTYlLhOpZL4bhO696bL2nXfPiVpt3euH7dkwfVl/l2ec0gxPgIfc
NYrhIh3426KyXF2h9vpAuc8Flb8sB+kEhbpQb5ARO37gESxDrUFsn3EPsLhOqz1o
dnIDwFRfhdACq2CTlbXE6xpdIG5KIA8lGG7MyMBhngDrPwzmSWKk6uAmYZqvbjll
GS6hDzjnm9vCD217br1xnH0St42xlwcjQUmgxfzT/L3gO0xFxojPqxX1dd+udDoN
Cknw1+cxzdcJ1/t292M5lWv9xsfSlc+O4ZBes8pkMip8w6dR3hVDXkO1UOFqj4on
i/4yeuI0MDmlvsg/AbiGfp0G5WRz+tYN7Ure0KX8JL+NH1frpJFPcWb4uCkIt+pQ
3WoP9QFrHODlsTAPG45o2GiiHNwr22f/rd7WoYYuqbT79ps9Yxd+xJGU2kDXUd7z
5Tq5xfhZVCpDpFT0W6lL8ZBB9rBIxBOBm2Y4KED3AUog4B/dr7auFCMpSBMVfuQw
Bq6kOX7sC3LAfolzrQQK0GY4W7OA3TzU+MCKkOJl/O5MkGSxoYQ8U6XurLrWzcg1
HAIg+Lj2b99n0oVX6oDYrvFsUg3k/NnIfYcR6hQSPWCj91rUhqjavQ+AFIRG/Uyh
+NWYD3YZLZSFBm9Rnh29WYcy+uK3kBQ6Mgb7JGC1jT+X1PhpC4obVMWcjdj3bQos
HaXukKoOw9MLp6DL8TbDTBuqC4gPrApSvkRZ1MGlAJMwvM/R0aBY9TgoT2CqA8uI
bVJ9IX6R74blDF3xzYRJkcU8WTXzv//zvxr0c1lCenOhzOtai8nkFUBT312wllbO
4khSvyZS9h3tOQN8+myrHow/5/Xb9NmKWRORhR9rkJ73tvQXr54g0q49YFmNDfi/
xo6vDMfA+0EMFHoNAv8oseM0zfp2xa1gIYJMlMRGsoFSiJR7jIIRcxpaqpErRire
h2fuIgL3SZ1TZB1uP4GCRJE80nazcrHbaarRCFAVepUVi6ffQPLFjhyp/aR9/9q5
MV17w+wEoWIv8PEuRv0CT5MmId5w2eM9M352R13ogvL/pU2cRwz7y7R5pH0hGEna
V9Q6P71K7XxSK1NjATmIShrB7I2bTx812635xbGRWUfVb9qN6u9ckmjdbq8VXTzt
PxhMo6pglzxKm4PRZqVPTMBgTORR07++7NlETqsFtApXE6Yvf6s8uFzPQs+4mEfg
2DEFHUrHMhdNGvS4lbzixXyw+GiyMAw8XY7XESxv8h+/m+t891CWtZQ1vhjJ06GE
GiE55mQwkh4sviqL5yL/VAx8oXANrarqGV16WZGaDsEznnzU6HIuaYRI/MyAspPz
tCImYys0i1WENsY1aiMersVY9sCtAaziCwhoAYvfhzN78b7NWuHtiDmzfrfc6As5
RsdIV0OJTckKlJnnoE+IidxOL8rBl4vKASHoGZ6soH0smIZS7akQxvySruatiXYQ
gGNIk2QbUbmGyhzmGv0oIm4cnpeTLyX+pdykosYmhbYq1sIvPlJityB1MnucIWCv
MDbpJz1IF1X1D62uVJ5Yn2a9p7nbdUg9qfVqi0N67IJxP0bVhx6f7KnZRWq3/mSg
+UeiqFxd5YQn0v6HTv0QItm2GOPhVo4xOpl4g8OvX2wenJJwalg26zxjL40BVKYF
zMf4cmHN3amY8W+6GAjujcg+Uz1vLElrQNsnfYToXBJi1Epgcoh81xnlS68pIlxs
yBpMdSrIdhuvXJVZOrn2OWnDr87ybQOTh8iqzJnOQjHvxwdDvo7kDYyryQ+vX5e8
6zmG7Qn9KmTomXVBP4g7UUcerIisVriRk29yDJxWFS3Gl1JLdFlHn1stZEEMJ1pm
j8pChWGMtdhFarr0oxLaMG5WPmQIiNyXCVPMHptzDTM2387K1vDRZqhx6NEbzk67
F4POF3Ep2l6hUIE18wo7jYSVX9tohCd6KdLMIiPu2NKrF/U4meGa/oYVe+gYhfQC
TqBRnAa4kpcGkdcOZ6pPo9zNM7ujuvzmF5JwT0fsZNxZZrOk/sFDsz8ZVQ6AeyKw
I+XIIst0grEY3ZlK+KAZMusVG3S9IhJkSxuDPJgyrTm2SVSmudXP01IbP/ITgQIx
mBjZnx8MY0pYXMWlwRQ5w1/jDek33M0bEQjKlu30MagVscsa6K3au+2U4g0JbzHh
IevfK2830pIXuWje8T2z2gZRjdpRnfgl52wq+7Z9ZvFyJJMPdTBOCMp/QEypR4AV
VCjoG5usI0tjMILOFR+ncTgCItetn9iG4pb9fgEwajLChJqb9nrYeHD82pnFvsDa
2082ei1QRy9UfWwooA7Wu2WyqJSkWKPpd2+H4aB/u5275F7/AIy4kDD5dHQU06Me
WqyO4CqpNfCGsteefOPJQVjIGx0PNLGwQz7kazmMJ75my64EoXNh65l4KM7Ble89
Zgo4p2H8t64Btsh9cYutAJDoUugQybbLdSQ/L3xy5XGgRZa2wezDr5mgYLaofP7r
5eUq9ZmSXjkma7IH7XNGRBbo+WljsUbs/fUe5biGnGuWEC1YbQh91U6RaHQpIsA/
iNGbRDZp2KjPUtETfxCGPBjxJ/+LgVVH2KJlAf4aNrig34l7QxmGdOyJTbxtpZ1s
mJhWgUxD+ns1OPOnIEMZxt4cNHoj/wGBEq0I9GjwO2y/UlUZ9GvCnH3M+YdcZveH
dWia1NjjK9nAe2pasky5V16C2MlJd8d/goEdMgPFbLjJg9Imqkx3CyVHaWkg3XWZ
SA3q7my01MTNa0Fnwa+ah9NcMN5qWUnFveNzxf4c+uPp+7swpRH4viJWileOsEg3
SrMdWa0UMR7C6juLIOB7JcE7gmCsDYBHNyoVITfeI2f0xvatj3teHT14+/EdmFRQ
BLjFZWUckwPproOUCdIjO1ZVSuxO2et4sevhweO+upMc/n4edDAIfaXtXEZn2if/
DhILw/A7g2er/11zgt8ufexi2fsXPXZDbaBFqrhT/LqC5szbnEcg3GTPU8hAdbQL
kmG+Q7ElEFjBFBI1AV+u/swwRex3ELAwPS8WvMrAyN3LU6JQkGLAYktRsTfM8YLd
NWhTyx41B/UEZ7e32KC+drXHGzKLLQbpVJ+0tdosiEeWQkuUxn6jqFqxdso4Kj6I
gxuRx4ZcGW7eAJ4YgnOG8YDTl7/528d4G65q1pMOjnK9yhkzIJoYhZmMGDLbF4De
nX1qi41ZHPM2L2CHVnd406VUHy5qPq74yTXWBF7PARq0JJHmCLqqNR8g9AkzcKVF
iKJfUaKcQcSP1gBAkLbl+zm559Vf0orhB2jY41hkHjeONa/V4xOvtmJZ97sI0YoF
Nm4Qlv3yBjeZLsrF+q93ZuvtPgAYtU8quhQ2zkDbGZPGLPdcmfItctDJb1H6avte
j55jVQgpyIjv7sQVPxKtc2SvvWmA3wlW2i9E8fTIRnmAs7tAfIW7O/VCli8QAFG2
RI6rOkh4ISegvuiR1X9EKGR90jxRgcWS7ulG/nKC/1+HRHoJmpANcf5Wj/5vLN3S
ugy9LfpXG3OH8dFZbo74DW8Ul5s1oltI5qXKVBGkOf4UF2FMED1/pNEbl48+xKIu
tbsKnwnuYyFtIeMMkIrT4eMQFpyuabpRrWbUxvYvTYZLAN9WVYYfy/ogZKOBKekG
2y1kZscWZ8OnSd7adN9cpWvLTDhOB1e0cWxROjPLbZJSlt9EzOLA5Abpnu+YWbMR
lwam9IW6OGRxZnOiS9Ph/3/ou/1fvtmdZsN5LnOvqkMA7Sfz6LXERYJ//dga5kuv
CXWFPMX/cKOnnhzbU1gwpxkDc2G1E48wZKSTKjT1HTCeggyefrVv3BRx0kh+A6+h
F9Tq/hW912isMrkm/iyrdxYGuSBuLHiHiUhE9gdZMm/F/jDardV7V63eY3z2K4xh
kHEcjd40TNajF+DsZ9NAYTfiaUZNv7nKLewHgKsmQvzuztb4wWYAp7OUAGlCrQpn
xP2IRjMsrVQUH6F4VXNs1sEfuKYAK3hc+GMrjR8/eHVeTQ+EEFJiriZJZ5bZooHW
FaGDJ6roJuNflQd16VvTqEU6gdIG693Xb1GwROt30rzrf1i68Clp1yh+ZUdggWon
ZWn5ZUEDd27o5yluGOqYO952gXonqmbJSnsGUUEladkWtGX2GsbsUqfElRCr2gfQ
AUun4ApobjVQhlEbuMJS+xfBeD4fk+RW9lhbS5TCDsxCBMpCY785hkfS2ZVNP254
zMMRsIqux+mWmGUbMl68dQEUkFMRRxNySxiTiY7u2wnj+FuNidGingcpurgxTO9+
FuL0a7Kd94HwGU4GI9aD5sA8qJxkQbKEDiqfb7csy/kp2styagOGU8gnMUm3uAOw
S6VRlHOFq9BL0Ww0L6a7dFgbeyJ/i8ic0lz8SUbteEhbAddqkFmHPbVX7r0npNzP
/yV7DX6MwVCfGAENeVlOnI8G3lGrA8gSgNktr5rquBm/pbI6K4ApnE9G7gr+gCWk
2CJCCMR+mPCkbjH6uO44uES2v5dB72uRzTpvAL8V4MOdYoCrshYDRHIzyuoCWShT
qa4PFosMaoZRso6OJvNf5HlI3lm9eG9+8xjqqTY5mp48+cFBelv1gzHt6tyPhW9j
uM0cQTGWbMPr3wwe+ZbpzeB3ZAQRYDN2tfh30IIWiyJoQ1Z4CeHwltsg14SDqoIA
YmAvdg8KmHFGfXUz4RP3T9IHMuzCAr7Oi0eXsT3ieT9WPQoTpSbzSnlz5117VNmj
RCVWhgm2WP+/RZCdfZvtkfRxJ2plKFb9KnW8oQEO80OcIL+kcRo4AhNIM0jYZbl9
/nJJ8LXAOEkh+Qv6BS1ssL0Yn+ZdPBMZt1zMoUQX7+B8Wm0vYBNMKGjswOF5G22K
6tVq1IJiWlP0jGv4PCd2RxI3/itECVJC2qtIG3be5VBvyDVJSKTz/TsmWYigfgz+
lSbGOXLu714RqJsOZDOdpkSK0HSdXORtOgW1DnBEiXo2q1kyh/dWhD+R5p0imLuA
fNoO2G+eIdGQuDSo2a3wOP60qxviftBz1kmd3RUdFbvGvvLVK+XQZU2wc+QynzDP
Lr4cQKr83kzam/OlKKHNcyc/U6beqEf7oYyLgNB9N7I4VcJIXe2Ei+0ht7zz/t21
dBQiXAKUpo6oq7uJBNa9iTKb3QqwGetoP3Mq4QpWjKFpu+yjQmlfwr6rnNRuGFRh
iD3BDgeSpq7L6f5bsbN0DLIi28T17AidIiGIpvS0ZInmeMobqHazWXfRa0DDRD8f
m7Djz/OsR1vkGcfRCbNTjGLkuafkB1XNtLhhxnL+jGCT++rgLf0SyXhyy8k3vxyk
VDIomqeiOSCRcp6cOyUQ9pJrun7Ae4PZoTkfaLAK4ywths/+ruAQC0nOTu60Ubtb
KX6NrTtp7TrXuNhN6X5v/WKK0E7byjAwc6Vo4lDW+DXPnTtJKCtBBgMxMD3TLAaw
y6rEiHAaHqLy0yZfPhs6JukT6aeZX+p640hNFYGWl8EM046gjqVMsnGe+QahDm2v
Xoct+WJfl7y8khnMf4g5DHiD947oLx6fRZ0EHYJNkasBnf4X8TZ85GftwLUe30JY
AJ3Pi+5xKLylTDdyPD8IeJ7zgH+Qln5Oxo0rU6Lzw5r2/NHq36SK9I67tWjSG3VD
faThuYMqWfttq8Thf9zfdV3fMJ3+eq+JpiUWqrG4cShOQkWf9CILB7y8cvJLhIhu
Q8dS76bGGOmpvNNxds3HwwBJ1NSuC20rJ4N53TBuDcDncgo7m9rJSt764Em6qbVE
aTxbAbdjQWPQ95Rq8K5lpht5TKzWnG/vmuVyRhph2l/2INa7M7rBD9WQNYY4g1V0
2hqVG/EJBDiourLiKEUlENm/PPgYMQm95h35HpY2WaCXiXg1LFcHUa6oOOGKcuTr
I1wVSbisUzRM7C0SQyPB29pXf0gEaiVjhJLmT8I4aTh40TujMRqZl5HZ+dcq5Cj+
6av+pA8y0ZRW5KNne4vk5OPsH9GFzVTutrENDzYHpraH4tMFdSjnmWPISMzraY4o
n4rWhA5O3maDXs3FqHVlhjcGJo9vjFw51Ugrc1Z5OODqj9GJY39461s9Y93xkdJD
lwtLGzoHbREXTSP7hNtCGe4EKXHDYZQIqFBhdVVu3nlO2vD5nGKAyQQxupvUjzh6
by6358gqG5SGdtc2O5aXf6USVLFoSBc9PftYNWDu76S5zdvMv4EO3IuULqmiGYys
gRTrPWfFqo+x6DbNj4R0f88NsBmPELLo4YZoV38MULvXv8+oVSypRHOX3Vi8oNpQ
rSp7RUTmto+8C4A9rY9XeOuCqBA210b7s2TUkept1dWeCXbIqoQFISiU56sCHRZ9
qOC/4o5b7JoY/uV85TKyDAYyN3u4OGjJeOz2cUF6uIlm6nhEaVoMwH4/C1fYjuVm
O7ftBP0Up5NbE/M1aMXTv75OY/xUk1jsd5XuvbRsINTOTnZrlFRxAwHj18KdLjhd
qJ2lDDPg8LHdcP+06fK2qSfKB7pJarwSqz9Cq1Iv+GDB5cD4khRnnkpVBTRgsyQ+
V0f+iG1guML/vIHuIhr5/Me6F6Ddt+OublFb3MCGQqe8wR0EQfrfl6g+Y+rKEZUM
yPrnfyAcg3Q5vTf5aYV0PPeoD4Obk1Nxy8vAZolxodkSJriZ2O0vgbDhJiLBF3MF
bchgN1HOo1bnql2Cue7cFKRMC3/PmtT+EiF7kJxfXL7Kb4RUStoqtDrY6bxuAGgC
2JHYFAqeQkdxDhu7R1VMgfI2OlLGiLbgKABFGLBD2QItnTKke34b8B7yQNAVo+ZK
mj1QTM/qrpNl+8IVB9EoX+PNADgJtSG5DUksnnhHjNgCzPo9TUo1VN09vm+WnxXF
iqRWVSsYwjL7vM1kH66w+LW/6yp0gOaJ5jZmbT3awOpezQkMRaUCrjEW5zcBMvtM
oFkUeXJgJYqrg5qFTwMmYF9Fk3dS5FjRmeTeaaFpf5LsihdDCK/QzaSIL4dT93Dq
zg6NPq5I5+lNhLHSgfjv6x2xc4A3li5d50X0UHmFRzU6thtNrsOw10uieOSkw8sk
FfUyV+zYbDF4P7e9S0k8GFLgmY2eJ7shF6bED5g6h4Pw9upmD+c8rNh9349B+7Ij
Wrvlu8RNlsfpPGUOtBC5YfRy199XbBdRlhEB3LPw69JOu48a1g4eos+V7z4ip0NI
oOlMDnSkzZybxRY2LbjyHgAjyHj85xLe/c/LxeDQpixgh9ZA5WGOpDmrSxu2rknd
Bd3g+kFhHbbBdF4yMxmmBeC6oaLTVwHcYztUZYMFo0EhW13tBbK/HLaZijrnYhAO
QBXT76dJxHntHkfe5G7xRosNtkLOyW6jTe3X8boX6dX+FA/7QHUFOcS0sXvapO6V
HOn4/3Bkv8P2rigcJZGhvk6GzXf1+t5bxlJ06bvToSPB3iNlNz8adGIEyaVQrq5h
Xe8Fm93NLXJ6/351eZKW4LfiQe8rip0c31v0PyNSbf0ZramMJxlRnPir1kFOG+DF
SLbmGs8qCFVWIKIdxneHaCYsj9NUwX1CyFIJ/FxXCoXMiZr2UJlGwDOUHtxMIXKa
V0jqrXNcq8/hSpnwP1g3tSjPlO72EnCtP3zTPqaOwmVJoPeIfHaMWJKRB/YYZ8TS
MGYAjW/XognsAlYclq6z3bzPKrwAR87sKYQvXbb5kklk96FvTjK5/7D2i7EbD6Ml
HNFgflgnSgG3kcsmgwd4xAgcxqS0LhU+n3tdJ9S0yPlsBqq75gPHJ5ER8Fp6hLp+
s/JB8S8SBfpa+LlQM4mBmcD5tXI3GhreYCIQ62lHPGu/ury8Ept/GFGL0mXj2OMm
U91hGb1OOMksoD1Zo8jpjeyjj0RYvLwmwpBjFepvDLty6uiSlemDprT1fHWBvR1C
ywLZ8hjwluBDXhQwYcjQC/8UZClQz8ZETsgZEeFAJKhzNFXSdmA1anDTb4U1TJ4s
LzFomsrs6ggtv7BdRgLo9ActAaorLwrAHUuGXIBMjZ5ws1hIE7oc/XT62yoyH/5e
tvJ66e5D39HqEmV8NAbk8crn4/htOlrpYAM12U+Rm88AV1T5YNR5aQW++KdPQJBx
hAVUVT30K1DSNb4X2smEyMq0BuPwsacGxRwCytUu7OUBNwGq88ONsoST62MFFuZM
NhBVwuZU2GuAXtqxdHUXHzKRROfO4yyqtFKP/jAbG+hf42VtdGhCJGyn+6MbAH2E
gYSnD+KnNliIyjl5JGRSfmw/pyM7moL7WqPpU5nFOe2NWah5ReZncUfGldJ/ln5A
Cr95fpmXPvSZcR77uFAZSX/xzBbzOdciyjkT2uYWjU7PPtC2hYosEN4oNr7vWjzc
ymJHSMiGo0HLK99m+rKbUEyeQV9re+uobSs3BxaInLiF6OspWYkxnyXGl2EKmwGM
KtNA7gZL95yTXQaKCkHVMDvnI2h2NIjB2BWzmPJtPe0ZLuOMmBZWwoTyj8XqGiHV
CTgrzzRgRqPe7DXrSbyPfpgSz+1k1246s6GSm9aSJTUBRNxKe/Aexi+QJVllXsXC
MsFaz5zIEc0ckA+3Dp8rj9IqijurlNkPEkWXHwSmh+rbCJAQQ7P0zOSFXj10iH2E
cuHiVqCkFwmnG7UT2z2kQb+Eb0pEm3ssNaXkqqzKLO4DDi/DUSnBbdS5KcGx+vxz
i5k2q8YbC3+wP5av/drJ1Q84/BYOy0UpQpY2ZuywgURIfMxiOuJ1ZRbCdhX3kK8b
tgXcxbLTf51FMWlSwH47GIRyyjETO64eNbo8I39DilMSv2SxJPL6cjWyY/pVmC+5
ZQNES7IG8asVmU+a6CBaH2ZWJgk14kFg/X1pNA/sO+DLm95jWKl4PySyXW3Q1mP2
OmBoYt9E8ANQ7i+J7hAh7f0rtO88s+87X3a8JxaJNXq46kEhXRiEZNB1K4G/QRxl
cCHqOE2rHrXi3SSJocFvSa30mAGilhbw/beyA68X8lG3GKGtwnkeiu4jzidgCaKc
rvnDSo9avs6bI3qCjlj5oQZZHATk0RVn3zDwmO98XoniD4XNmjzM9Kztxl1zHLLe
rm+O7ApnU/xYvqp8mqNoq4pLDnoPTLsTzc2XIH8gkKgM5fwpN89+T8vvZp+GedOz
+yeQalBwQjpY6HgeOlwpjnQ1muxvvO3da3EIJcmNQc59tt1/ZjuoDybbNUxrgasQ
izd2a7KdEJSvF5cmf84Xc8rfyWwbYkKz1ofu20sgGg53GAuAcj16tRVZe51cu8Hq
84Uh1zNGnMdd7OsmHAwL0nU2tefq3zOAHYoGlOgFIvT9QFkvohVJPQWSrv9kzX1Y
obVaHrS+paZ2uyxI+a30lX/x+Io7c0C7SzYk7LzmnPbXDxjaKQu6JL7Vr/1114Q+
eg9a9osjwDRoe5uoO9jzkwD1yKz9krsjf/eUxgMufea2N02mZUVUgITUxW4b+Pkw
1nRtUn4UCsz0z4TFwYSLhWEHDZShn8vCDTg2Xs3uadqFjwiIfzrbWlrThD5xQ5Pf
3sZxV+/CEy7Ywv7HuYahCG1Ae+fzfkfS0MAOndsMVF3ow39wsS/W+h5tn9/ezXD8
QaAnS7cNmwTHLngej1yEKNUwqGMtRKB7CAhcAh42DPXXxBbuhzVDRDHLcii6tw2B
IZ/L5SIl5mjc0dD4g96U43ayVBVqnc+fTO+EH6Akq5Ipe/199oN4s3qXiPErKTQQ
OUN5x/v+o6gZr2zDP8pvaKLl1DHus0LuyqGjCgzEFqeBnYXyNXUD5pTIjbYfIelP
4QhZIQJVlPW4u3ogWEr5eEtleCQdvIXs1HT6rdIenCRvsYWcoSJlMf4xqZnOeIP6
3fWB/5qNJ7Q7HfUmyiKpAPwZ8i1n3+DaovPICj6bdjnAbh6E8OM+AxYQdYx1P7Zy
O3ZAxqKtEBElAjpqxhSNYKNiRIE1RImIHGMuQY6FA0fOLMn8iteSyik83fpRgo2o
lxJqsMZ4o6wJbgsff1dEW9BeAwxUCNL98rOsOZL1YflLCThYbpMX3t++p3fzMwEd
ZMY+4d1UKHb4XLkg7CHmxs0d7V/00v8Cf3IXW+4BbmQ8ETh7cwy5iDmO82y0VwCJ
Hav+8Uk/QHfnhQyTCw1NScg74AM3zwl8RM7WYJ4KsiHmZs2DGMwjFpIKV5Fjlxdr
OGl1kernthQlgZJYT55fqHNeDSO5GTeFCt9MyDjey2Q7TBTGZ3eh3+DVY4wZlkU1
NN4bzWJBZ7wg2vqDikikW5jdeL9jZz3UjUn6cXbCWdyjPq493LyBYYQK0KrozBjz
bl4O+UzfWfR0tRbUEv72mkGM/J3LdY7akCLuV0PmC96HilUnvKNhyE/QwAAoDJMy
yWo2X3rp4mgPggHoFQppW4e/SDe/5BAja4PqYgFunYHu8jhNtWvjKMwVLMnFP2O/
EEnYrQVOLSi8LbeomCDdr9wCbniTJn7XmyJdBDBSYXdY+2OiZEfaQA4jMClnX71k
qX7fx/4VtmLOHck1w3CPh5XFB02xu2kf0y32Zdytk504wt3yU17UOEhD6XKVkye6
0BhE2v5cPY9fz8nsA1KFMF6qZTZgZsV19jkHia2qK8ZABZkLBW4vQq2/pf+t0bOX
YRfsQYzabPGl6nYqW9O2AXk5Asicd9SbJb9eblIlUJ59e8Bzf0+dtsowg85plVlK
wdsY7OqAQHvBfWu/l3yCjv1J6fyCCT6N8UVtpUy6+jmQjpBU2/dthrbzO/FY/A/v
I5Y97AhJH906uHATKlUGuFBGmKMq5EQ4RgmPXZysGOAmrBgGk+sl1QnlpIeWSQlh
ckmNRWeb9wFOs5em2dtVWaE+A5jANFn5Sfzp/z6cEiOM4LfZI6jwvV/dWeKbjENo
NJBFrgDyx0pUKWlc90eok7NSOgzdK9Gq9EbIw7+sYH3ZSpklr5kue99K3CvIuEL7
M5x2/nLmEsI7vsC2zBioYMnWkjGCcIgR0s9OKW3l7Q5+uUjiCB22YOjQU5q7qL8K
Jva+DKWjNWeJ9iHSos0JnhIAMJFDtzAhuCCwonSBDd5pHbGPl1W1whWEKGmd+9uw
nCDN7hx9B+tr6P8mQaqZQpJhQNwe3IcjAk20y9jtqCd82hx+SigLgoXJE87MT84t
AjFH8W19sK+lW2+KG6KM5YEQzeIA8p4ashkzQfjBE7vn72/mv4roQRh//0Xx5n64
ujplAbZeWb4FB1Z1RYgf7QksAtyUFnnCUA3L1CMijRgbxr0yTC4/BO0NbKuXy+R7
ocf/N93FIBn1lDbHhSogoMJOPHMvNOOIl1icmLmGmmjDw/sBp2TxgyJ24CMBy735
iQ0/t8vPQefKvwMpotAAI9g8ZLZEMHVZOLUlQPI23QemknnYTwattd49hNztkhf5
uw2N1xJd1HaVAuAkOPQARb7iaF81MoFrI51S9bCtVMnAM4c61/UZzLJDJ/Z6Jpyx
NOC7hfrzXTIsA420RB5eTUSyrXuwgKA6jaP2kflRqW/4LbHG83J070afuy1wzcH0
SHhl/sYaus5lORxLHH3E6iZcVgLWy8KhJSrfTm/LZ3L2j2aDzu1TY+573zqyB73O
daiV72ifqDrypxJLFR5vylei22C3fMNMmVQRZBF6zOQ3dQ91QDJvnzkLh/e1tLkh
rZrg44dThfydoV3J+nMysBAG6uZL13tTK4/eYkzbNbcSrZoSx+wMW270H2thgRSW
RNJV9b7ezfdZKhNb0JZeNUsfLNE0/WzY8CcFyC8XODJFsxlcTSnKmqmHieAS6Gb5
x7W8LwAJRPn8FnYFm/luZx+KqAhBP/FMyeAsKj7TZnGznAs76CYOV4pSR2U50rev
mV8WWlPg5ytN6m89JqZxdS3rlxnq+fdeA9UClqusKbgs7R5fEsMg7D3CgQS8Peas
nJqu933K+PAefHymPmtkF0YC9lWVbB/DLCIaf7NhndZH2eUfy2kC/rViE0sebAZq
dgc/JdpF9FuRyuH8QmmiRKpnLCRwdcB7+xbrk/PtsG8oqQP2IHlnC7B8dOBmQ91J
EiO76CszPAPluLZr8ATjpnUAhJJrNLKn+bFUDBvE91KeqoZO3mKBuILoqt+ILRfj
i+94In/46n2UApRzJnKnS2Ohg8rgC+OV8RcANCOv5TUuLczF2u8e/ID9i3Lv4Hvz
C1tfch/R4/DtrcT2qk77y/LWhHHd3sjVDtexx6sTAcf0teMdKiqnGvuiBWs98oQw
oqAs00U3gmJOjsjA8FHfzFUOI4mK6qXxyFH6lyHDf7sEP/BPeQdMAbbv/Rbr8yco
wsgQoYGwsUuzUEDp5kvYBaQO8teovHFT9BwlzdwvbUCAzxCStXo9PyhL4kg3a2yd
vCT1KHwWIKFa2WR/Ku7YZORMKcUoXUh+dCdEWkD1FM6A+91Tf23gtq1zmyE3NVwS
3x3XIyXCn+dtTRwlvu37Yi/X/mgI3gV1MbmNRILJ1m0iAgfQSbMKt0JEHnYj02iS
9E/nvOgzR+ykXzZyIn1kJAQVy0GwjAM4jPS6e18bkfxieD6wmzOvAezVQPuODqiU
U6SHvAjnq45vsPwQ6EGVZJjvirm4bCVMiooeMct9/mGBhiqwswpfD8QA3GVNFx1+
zaAFZFuWp0D0KCMKBP8jONaKp/ZT2SYHSu9D9nYgjDm5TtJOLRn3cbBRGuU7a2ic
VzjjQMKy4IEehx+LkHYKw5b8Wqfbe5EGNOCBaeeH9l/ICSQCYGbDBmYWXudOptGD
ve7jZn2iyhmKyzYQigm5yaBeZEF0cu3GLZ4KyXc299gjoxTyYwxQq7CYQFWOksy/
kRx97n2TYqV1iHDbP+Ne/cmZIA4scqeivGU1udwe1vzL7p2WkaBiz5sMxj8dd2o3
Q1YRuerMFki/abDFcoAj9PTWIV08B5ETL781xz9qkxJaSziHr1LIBtnwBML+2b6z
t10vEpo5LQBF3gsbKjyYpR3PemPUFO3lnPETT9sNlcNqE/fr9nlaOwTRv/1EjrGo
zMVYpzVb2JsIiyn09CIAuDLYts7S17gNDPLtTItkfkVpAHjuwAWR/Dvwx00r7ipw
lAyTvy6voSKSVn2RaHuXgXjRnmHj7GtX0/7ZT5mR35+eVXEYUnZ4qU6IqAOESjGo
1O+jDhrpZKoJxULgaHInCz8VuLC5tKTjn94EF42gUYpzxIrSMm175ZC8y/NWzWKx
X9q48OdY3qqaQ7qNw41BtoTOHx0ucRDd4gVNhn+aAHHmoA79G+AwVTQK8TSTrOyP
n0j8nGz7M1FArdn2143nP2evn/RmAQW07YBzXQo3qmGgC5l6dnGIq/nw55hx5Fvj
l0a3rTx9L7i7INceKdtI+dStlLd63CWxloSW2bTAWmkDe75E+p3KfaWwicZCt4Cb
IYhWYPDU2xrJkDbGhj0uB0rlA9uiTbsLferMpK3NWd4yNS6Ei+RAkE7FUW4ylKWo
66XcQdNO4ONbmR6/C7F2FWnYSdo2yQgGTM7Vi2Evtfq0k/e7S4QXHrLU1AWfUNaK
2SOZPzN0jjUv/SXW0s1rNJ3rANFLKGuWwEbudw2iNAaEnJQjO6ecfApYn1Utld6U
i6fSNb9/UJSjT45wdVI6ZjS1LkiDoCn2P49f/H49ybNeigYES8xMGVTjDdlMTrjm
Dd8g5plSRjdADBBnCqVMVwFlF8JWc6FwOyCaEbzPN5NXFsTaNI90x3ZjUrLo1yTw
cR4dmzLR1CULm4sd6ErE5R98ncRSPD3SfwW9xWzrUaqIZqEJm4qMPyyqDWlI8A+M
lzV/F1UTq8UJSl701xdFf0FaRk8aUcD6nNm5WxLCk+xsDrNX/q+/eUVy6igC3gPe
BxZvKBMJYoy4AcQgDIO/F+Q6YLjQ0ywg8dY3N46DHQZlby1xZxRX4y4oiXB/T2XH
E4IdBvh1hsC8QPkQMN6Yo/2l569taWJxPpauNJNQA1T9y5vKk/48wgyf9IDOm4jv
KhP50Y1CZtzhaqiOoFhe/0ePUNPGOpB8GZ68hXPx0cdENRIlA+Ke24GhNskeG9fF
8y49k/Wt0+rYK6mPceP1x26pE8qbyaMwA1ZhhZ2Pily4UTarWTa/SPZEtA55FI/0
xCURRR7VHr3YcwzyOzDuhUJvX2oLRFzzAH94qofnGSe7SBdY2Bnt6192obMsi1mi
ony3s1DrwzSIB51ddeBOb+/AMyFen5gkbc2DzH7wVoanLeXtdzfLjZ7AIO+dbpA8
YtfWFRF1+3XgZqWp29b+PjeF+GeTeEdvjp7th1glIWDOWPXSjY5r9cILtFy2XYmd
7E+8FvZaeQeB4FZBFNaRXyvfNi+CRzKcH6R1YgbPdPuPMc2qRKJLIToVOPSwrqzj
JcJB4IUJZ7Vbm7zX1T6TPqyTrN0NdOum3MBfozfoMljULRQf+h41h3lgzzFlVhRb
gZWcaswlR0Icg1eapjRzxvbIBhdr+4DVMKpYIdt3V0OSumtvUX07LVpmpSjgG3sA
+hX9H1Kiri+qAUMdJgPAQdK151enD5dbMZ2izHubkjHJZvnk7JGjEGSkUaO4z8Ws
HQQr/DVlxzdLgxh8awOGEvIgMBTjv53C2WQ+NLNLS8oj4dhsQCUOv9jKouu6B+up
mMQQrIZr/5Yfv93iTU5OgIhvJk2H/nJRL02MKyEnPEWesrc2YE/pEPWhD3qQEDxw
kfkJZxBLJhdrUMQr3j8qsP3cXzfNIxHoQMETHDZL8EwTIuntuSZZywo4cEkifJsf
DT1fZOxuxTdOlAb+DL3nN0iFd+QVApTtjDVYZNFEeW/uqyJSfVpYN8uFhva9UI+a
YQMNCwzjwGFXApaa6LOru+ZQTbuCefO/5cyinVfnkQaUc2vWQ/8hAVhLTb7HpsL0
+MkjkXauvRBWJiu/BexmmxQgk5M3s2rboM2PZySPO2mZaiUu9cWCyK3yP190Eto8
vk0jkGldystoQgQX2zoIxvsv56XOjLDFner1jMCR23PsRHRSRRm3SIPkJL7Ea++v
RO8qLbEuTdW4arJmwjKhgicaI3jhnYwDMhH3DwPNTiY3NIZ6Dg9BlaUSgb7XszDk
UvlB9P7dBQBETI81E3ork6+6bcJ+uf7O/CJQU2yWvz1bQdla3jEWLxjJN5m+Gy4D
Hp5LhoKhiaxzyrOxZAxvDlrwX/qakpqujikxv6YdShh3R2WJnc8kREGHwC6enOxJ
BqpCK/VikEhGvT0wZ2W7Z7c7Qn4eTvAI3bWpx1uiM606M+hcL/5dhrQKyS/EL+oS
x/CHU0pr6yIrr62ZxTVSa987RAC53LpTY8h+LpK57c4kcPjxgsE0Oy5VqaQg6c7N
Ewi0ha/lJrrX7nE3nTbUPjeRUIJ54KU2JB9jWuZBXx/Nr+s8/iPa7JedFdY1lGNw
mVcpEk4E32rJHXn9Y8o9mk9XuJAGV4Iy/M+mkW/hnof92JzrlbKI5hszLPrLXiVA
4nyRAMopMwIdwL1t+b1UEE72Z3+ztuPFcMvLXx7YBrYraoPJft+Mwfe9YJPhgPOw
EtolnrmuEj8o98mCuWxgFilUIjwK56x//GU8m4CpdoyvYvh6cv+qZ9EZ7/wlm+AM
3iSmywbfC1hrH7Z/dJSDlwsrKqQ9zru8ZFjL3aA3F17vmIkZL+CKQl5AlwNbbY3f
gCJ9aFhXAAeoGrk3cbPaRKbbnWJ2du7zP820ECTHqwOjV9YVjRIbdhMvbCLAf7RM
DAhNUEs9V3lpRCuvRDsv+MyTuli9rA/AayGJGLrqPUX41bfVTfbOqCMY92IDL/bS
/UoM+cPwHNSa0HhPAaSY3JpsleB6otPfe1fnvcJAUTnEaKRddyxaSlHuHQz/HqIl
LatjRaSWL8R1ydpsluAXnoBEkecdUglbUDZNxxjq3wUrcFRfC7GrPSI6hpK/yc2N
mlGe1QF8b9ynziEkOkpLlSK7UrfHjeuLLnr2UvDzv5U8nOQTD+SFIMYFwJBdyPMw
EpUh2xhpe49eQqrZF6gEvEomwPkiyT7O3ZgSdIL6/ge0RxluX+yLWb3BgpO0FVi9
A6ndzIVTcxwk8UkrcVxShqzAer/7ZEWK8nUEPMVcDC72ClRo8+M1y/FXhFx1Ycao
Zu50Pit+shYiherRlLAMCS70voPX/LMgGyxt9oe+eZAbZewhdximYJNG61vjJE4l
YsR8sx7F2cpl2QxnoF+9L0ePShaFTBsgDkACDqobsbFQjjbtoRtRA2eUZDTHL/SS
fw4IvpfY1iSTuv6bTHhpjzFzMziel8Pi7FvordpFYB4ENnzg+ESp3BrJElOt746+
hlEAodxnXoPyHBpKGMrn7IrfYI/kcpAZyQQnFFM9nlrOdsCtj+nrkIKt8T5r0akZ
iiRZRAOoBlgmqBv9lD2VHe4CNspYFAD6DxG3VxwyjykLKdEZ3R7Kwp4+wWT6U9Xw
yL+GomYJVpT7SEZ3PB8BTkd3Eyn4//wxhxAdMrf/EvAnM1LuMIK421mM4e1VoCnz
pdxS0/r9LJqqPHAz6w+69oYTwFzzKpmNwFO45dQDC64hBNpxELObw8cnI0Y2IvVf
pZN/2WHLSNCdcmgeUpv3l05nO8gktN7JqJcFBKg9XOAmFuAODZGQO0AfzfemQIdI
I8pmk9yc69CnFYzSKmIiKDabFebKnmNYaRst8/S6y9aBfRbK+e2Wx+Ou1sh+mkEx
5Yws3J27/wl7u9fL6H0unzW0Blpmt12FZr9rGnpmgx1zXmJut6QTtwHhL+JidkCv
U3P4IiqRYzfNOb+emD82r4CTaAlP42bZWokBaYeDI5Tim5eRjwVN562XMartOXl7
F8rGHo6tC/Jywx4zwU0/4Rs5DMcEdD8bglo0XXG+Vzm4tMxSW7fhcyXh5/8WOpPH
dHDongO3VMT5a1KpaPl7zCrQnQpthYBvtxPuxvB0VaegB0UN5+KzxHBIM4Z1VQpI
ePJc+a5S4zZ4L5HcnIO+zsrqc554zoo6p6hWXeLZXEmHwyo/ihyAB/T6SWXGz8qI
3waWr1wJciXGTJyJjnH4zs7Q57HLYVZEvWnLS9kBZYMzB/KER7PSR0NhL0ihWP5F
k5eWYmKxuzXG+1CJMm3sGpZQvNveXwLljAunRlsQfOt02Rea5tXI2UNH2Eig/yQb
4c8YfGxNOPGJeUDsmJNltylkj3DyVby17gmJohBr8vwXI05gRozfxswBWuJ09mbV
qkmm8Su7wf5xzAD/DDJ6OXRBo+6QnKwjcDYvk8CPPWWW4pOZtvFTtD0JmFFZtZts
Q7PBzJw7/qxK3MX83TWgPyXlS7VhP/08ia1ZBPcv5KpOI9gftrj3YCKkb16rTSYi
Ps9eu+lAlgz07tIE3YNufU5bEvVH4lX+VXNMVQPgqyC5Lcr8l8WwcnY7jft/bV3s
opfkt6pc1ZUzFt0mnIX0EmIWStpoRrx74W3JuE+6lg8fS+IOstmYsQG/oLJtP+6T
gPPNB49gRY0vNHI4IyHyzSSBXQUeVOFTaMI2ZxhoImMwCNfR0gCcTgLwIGHUcmZj
244di50vwsmZpMSFlC9Ljv34yppLvY/uHJV07Gf/X1juDZyggch4FTJ9RFS8SlAN
fzlILoKFjLrpCK+uBs+tqwmL5cTXmih6Zfv/n4UnIvs7w+tRXqbWX/q1mDGxpGCt
lqTVOvOB2Vwyr2A8TGEjW+1H4Lf6vpVdPwCRxhD0HvLz3M7d+QxxnixToPVyHYZH
QRVyBNb8LNtj7FoHCuVxxZvVBoKUi7oc+hg7GXMgsRP3pQoEdhB+c8AkWdgu8ugR
IbpJm8TFhY6bvYounvNhCIiWSS2VgwWXnlYKK6nOmcNn6ixAF2/LpUe3ocS/kCsE
FjaCSQbjva/3vt+dNRg+lIgBbQRn/saUgzCBuSb8RqDTPzwMTy+4DNdJ0v7HjZDk
s8gzBG6T5/QxO6TCFFKuXDsIZwCI5Ok6vRVE0sOWJ3QhXJZkVmBxBriSyrYVt1wV
6MCVxg7rrI0RmKmvT40QvwvpADvhDsWAopqQq6Y4zGZfiif13q0PBe6lnFSb9G3H
nXTa6gcihwN8tXRuX0nRF7c1psnTTwO0iOe3UfY02Kp6Z+/wbdQQv1c/+yAVFlfK
/P7sSmvVZL/KKBraMqvX9+osNOYf4c3cosblW2nQ5nqhBifxccAxj9kFu9NZrnmW
hCEqAnNNCwweuKCM6cuxPgfm71Rsf8RcH/LiryEm4Bzx9H5Viip9r3r8K3XMZX4/
AeOopzrlHVqpfOvKgjQulL4Q4SVCd1V7d3KQs7ZZb8t/+v6WKF5et34YRlN4HI4p
kT+wQMlutdZxkz/agAeZre0C9mVLXZQLfpe9FW8dgfR6YFgUL6aSfq+8Yb7CZypD
Qro6S5/JJ8pAqjFkJrCLAr3zAl7Cqg5ZqwUyWhUsZPL20J8WKjsRNk8L80bnpI7n
Qr4uTVYYOzUx3iYOZWYBGtqT4KArL1LHJ5WhCUimwPWfuXiqn61+QzSvNSUZFbcz
Ifvn3BZlwPpF5MIgLD2GuqfzAmLA8wtwHkacNahN9oc4MvYrWvENayITZaUUSUBA
LfLHSqObz251/HZgOt+e3mpr+x9dOZXPtDrtOsR2HUx1phvfOM6diwgBFOdEEUAO
42mMI7DnAYLr4m+vOETuRP3YhB4pk/WZ9TKf6QfhibYQTAywKFVKwzSFt6nQERLp
pVKox8RqURw6psEH1GrMXOzk7gyOhY99tjTXNioVrgUFeeIaLYSyp7KryR0yBeBX
LOahOhJUS8kXmUN5VDpBw6EGvRgDeDYw1HBDHGSotggtV40XdMSqkERSN58LAjRc
7PQOVizdY4SVcftHHAn8kqESNv5iPGNqhy7gx+OB552mhP7K5ime4U1+nHg6rDHm
Jh9AzwcdXjVg+6tGOEZVg9PD1zrLdCquR+UI1Ol0w1hK7nnOmYIH1hTcILXQC02a
eHXVZJKtykg+25DG/ZjCk1fVmnId43W3gpw/OQ0UyrEttXmFx24C3HivLu9hoAby
xIK4/bYD7+40uD+ctzwACJ5LQx8J9ON3xeJzIOPYY3XKzUpFmANHhIqpZyVNuHci
wOjnT9Rn2tpiHhuYim4n33WjCmRuSqHaydMXQF5XDLuOQnuH/OfFZuSznHgujFc5
e7tkduCurCjZCUbqf4CC7YEFWhTzwE3RpRtxQV859PD/RWSUv26xYNai8kzgTgp6
QdC+qaAtSp2vn0ASoz5yTZnQr3QEiz+X0LtbzFjrHHuCgKg6TJ7YjD1M9/bnShoy
Om3MH0sZwLLb++Fw25420EDViSrJSQv9mLAiKmb9sEuGS7Px36yIdZCJWspV3cne
gOLK6bOVMHVpAWFCKLacpkWcH/XxNPdIQRAc6346YD3ZmFwIsMsfsoOME9eMBXWz
5TOZze3OZuUwMr5/X7Rhn+06jjMhje1osCbXo3dXtyipZqZ9XGi7TKAGLEfcC08/
sfSyJSc40WcSXWurVjDJQJw8FELeMIJSXQU4ZfMdKaFQOsCzJJV9PwdpTveVBxcr
7hGBjiyoT6GHAH9yCNHQbxfZHkByFG4ZhsI2Ai5yko+yAkLm4+su1wUIuvFJ0XuI
aPGOD1drVmmfYU0yXElGc90j18Yy3rIR4bbsAQTcNMVXar4Cjw+MmEFTYZlClkaC
qG7+pzVWq2Km8aT4L958Gv9UXa5COhiRRKpYZo3e5FRjzknJvmu3c9nNKQl8VINP
9Vp/UbKUeW/DG8ZAoza4TBILcpsbG0S2fw8hOKr2ToVIXQYhejDx3w+z/EUmeMvi
0qM9ZkbM80+L8WWjgzNFDWd9Jf1q22oZ1pcon2K9F5uVg16cbnjegjTKg1y5Go2B
YPOk8/7yUEip+xpia5lNGA==
//pragma protect end_data_block
//pragma protect digest_block
7P9Y2NluALNKdFPOuNKpu7+659Y=
//pragma protect end_digest_block
//pragma protect end_protected
