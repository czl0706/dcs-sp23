//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
LB78QLw1kyBcSZ8qWQKA1PMpzVzEuUjkuwJK0VuzLYesD1sN3TZ/gdH4ooN5cWhR
RE9zQ4wdYcZl3Kyipco4k19wUoBmlvIQ3azWPG3MU4sicU0N4j/LHDHFvmtKBWkj
1sT3c/L9z0pn4oIZ0GWT6VygRyM1a7Q60gwlKW4pJK1OFoydcrUbFWatlGCJwRbM
5XiN9+wByZl8MIOdDy8CMv9/l5blzzVj8QJCnwWcK1Pc7rRFewdiaqxAxAokDRV6
oN8DVAzyCZCzAE3wKfERQX3LC0cLfIPkjeT5t6s1a3n+Ysc/kkQoXTKuDSotWuGF
p0KV7h2Oy6mrT/X2R75HfA==
//pragma protect end_key_block
//pragma protect digest_block
pDmJu6mMoBbrQARlY3jV7u/3x9k=
//pragma protect end_digest_block
//pragma protect data_block
V2U/OGv900xO8kxoRQBRVstFiq2OTHbG1IvFLUxBsx1lcEq/DmvOgfNy8HZfSq3B
tb+erUp3VlGgXvKbqDFbcZHOsEfqgFzfON4hH/8QwDHAySSnS7NeAUNvwvGadeXe
QeBaKiwX3elIzerHucJgpKnkUPTQOCNYJAxeY3vyZj2mF4npeC72xMaI9tA8KTY9
Fe5ZpoZmKneX0xhnhynTM1QolKB+n8TbUGQFeNj79pJBiwJwdrpYCV6OkdgQF2aN
5gdGRXp2FA0k/5Pw1ltlgz5wmalXpmyKuDMhMCw2Ml2RPEEepiBGkBPM5xQG4O2b
gr9sLw2WwE7xwHYTPU4+is5+pyWWdPx6T+oz+PQnjc6gi6XC1rbczJAngGzdSYS0
WKecf80ddmbP+N59CzsExHrFsLLK62n8809VhFQY6q/eBcyc9Q2GEwJnD9j292wG
sWdjjfI/7JpgNP3IwohQVbfMqlGDmTLZOahbG/esjMfSVzU3JB4nAWq1B090NbQi
xRUl9El9p9m1zJAUdJOFA3CkRmCjL57lY1qAgelGBS5QdbHKipVrIA3NPCZPTmlF
Fpy/k9qpQmOwvZGhq5UEyWkvzuheuc6xsyDXunxYhpzmxgRMBujZC6APO2lMzzSO
Vr8zvqMmiNsY73IIB2j+6577zIvU7Rb8SIgzmOKXz3BIo+lOEi8GEvWJ3TxSTeN6
NejZ9o6CsulCd1tK0PWbwM+/6o8idQo5CGTBDWCy3B/5DQ+qzlvSMK0v/GnoR7vY
K9EPrrT2F/bi2B7mG+Rk6IR9H9Cdg3l1j5+aBYLwFv3tjJpvBzz1UjSm0PhcJXO+
CEFECdQVhvkWQYttIKp9GzmiNCqDLcveiVjAXxyVF0GkcK1aGy+40CH4k1XOT6t0
jYLh7e6jhKx+thVvUPgsacfzCJHhS1hXfIgNZp2/5OzHIicOINijKAJ2H7o7foNS
O1erKc98vvVG0EL3mIMczAf3QPaQ+3W2v9YUqKeMHGAkNOjEOyscRwGTjqeqp/A+
x8UFQaO5qkpatcPUAR5pGIaz2e94LJckKdFHIlNumTarfFnNkcQjh1REK+yFCtMm
nnu7M/KX84/GVRizjYKmo554mpyT3SuJl+HHdhTQ4ua6gfsW/OqRXHtHFNGi6bio
cCix2Vh7zFHkiPy/VOdD5MgPEJyyRuQ5j4o/gOeg7tkDMUQk8FGEaHuOUoholykZ
3o1csPvowkaqA8fFiJ4I5ZYXz/nLIDwh1vcD59+Ffy70lLgfPwKBkoRWqA04oMLY
Cl9Exu1i2EhPRqSBwt2mUjJm5PBzCgxHPfsYWhM7FagoaUUuF96m2NHSNzgAP7Sk
etpPnmscs/Q0a+TCQo63DgnJztfcyTmtWXv6eSaTpPmQD8yQcvpm5chxruL7JZui
0bHSueRjo+7uGb+Ai28qy97u/af5l2ZqW/feYv4UB38KLpgfhyzbh0wXtQqSWOeL
PFhow4auBzJ7YarQkihxUatRgaGEdvZv5Kdy0w62/RxyZniYyg0WPsmHxZpo6Tn9
kCHlIz+68eDDStBMsRfDLIOHlLEjCQPvGs8gfCscYG30GEGp0RX4+BWHh1s3ENfK
DM+uZelJirYSJgrYa0ZbM2DbHj/Q96CSl9MU0ssFoJ6D2ouVZQrlDWrjHwahajdp
2Gx8n/XdH0EeUj8cD+0TyUM4dqQ9ohoMvOCPMcxGjIn1H1TXkM8ZUoKI2T8T8tOG
axIJhoE2VpLZdaABemB+kjSmb8LN7bbmp8qEF231NGiU7bP2StfTZ9OnK5UMXHBY
Xzqr2k+kCFK2pTzFSxUSz350jvXqFfHeD2tp8dzdT5Jdp8XgHgubRny/Rjymxa+o
0hmoTMtLymN31GhZWMUgk6+tlarYVVjAwD1t2V340vl3F1Y13xcoJ3xE+MmZKEyq
Bu6rJNazLSrRcj/p8p049i7m7zjJEOtpFj/AMBZQtlibRBJC87FUVm4YS1grh8n4
aboiGSFYuvEfBNpU6dZsXsQsBXwi8mE88ajVP16zG3cZfiC+mjdISLRebc4NII4G
Evywkj/DedYGfTG0oCxaHY4eIS7ecciolXuC9zKh2lKRIZaw0dY9sTJISUAGhMJh
a0txzAzBnHa/YnpR31tz9nXvScaaWLInXZ0MjY0t3GfOzxUVfgUhxFAIS4qdNP/h
go6YmxVoAKlVxcvVXhC4y0mEPh9tMBypyHhX0DebZTb4eDXHB19dNWDN3xYUxy4V
2GuSgoIFH7vr9UQJiIFiF/9yBmLW03wS7cUrSrL/PYzBHUNsZ52aJHKbwQf3G46a
DFiMjCNMNiFLFuOCqsXAKUF9ylhob8aOd4Wc0hnwse8RDGj+uIz4k8nSK9cD+CKj
HKj7zPftpbgF+DqhUcNvhIHTO27rKUPMfH+PKxDuSyREEdHfFDewMDF8QLvG2C83
NzHzmweFwHis5iaMAXwCtqefZsHhr8OrCEPH67eKWeofDwZdZz3nJTUp0nT/sbnO
lcnVgVfzIMAgL+OplKZOSqZWUWFzB8BBkjQdZT2MOjVWUSuXgA6Qpt7uZUReA9Pc
lHo0vMZxU3jMV8br5hIsb6mq3pMqB1rT/LYQE3d3bd29+AQ53/+31J88Ankg5mjr
5nhmC3gDKU+baWZMIuL3Kh3L7ClCGK7SgdN4/mUtcX9NFW5ZuWrgFz/DuEptXnlx
0Xe5KHvI/xKKM0jhZ0avwbRDjskQy77ymaJeGRqQj0ADDWfO5ex7urz565avRl1A
WeAbo0yuInzekAFUzOHdICYwe+VInR0gFSOhkf9Q1YCis04GtAYLV+B+B7dE07dl
Unink/6mWZi//XnsuYWV8T5pGOtN2tf9dQ0HJEbWBl6kuEHh1GkZAlt9yW7TlorP
9spdNgr5hduolxdzEpe/yESTaphxfaNiyKYwD6j/n0tZzuVOepfAxuyL+knxuFDL
FBYAOt9pzlgt8uHA8SU8W5Z82BaLoE+sVb3sfZFxpe8FQBtrqQHQW6OX7SfxKpv3
yPMvr+Z+gQWH8BfPSBDolAlWX9d3vSMbljDuwwRBeGdjMfKdM1nFuF2nLU/eeDXq
Anlp1RcRpGvnrcq6Bj8+kn1KhY67sDZWRQm+mw+fsQ9+BGcoX1Bv3hs9wkdn5Tt8
5vy3fQoEj3zoaFsQQRVUUL+itQwnCkRk4cZ0zWitfntjbuWNfNbDFEELQCD+8U3j
fU7KMbaCgW33ZH0eB7YLzYTRO7J+QXeC4DpvMMc4Osb7ZJW7sg21TxxVmgWtVukI
gpLX6lou7mFBk2CBRR1EZxnpaRiRUuW5PkkyvUONV14oqnls+eEzcwtG9GXyEExt
O5moH21S/RhP+eYa+Mv9s0QSKAHi/t98JKAnsDhuFD9n+r3XZ94INj3MxX5bbnGz
XJEFx5VCXlfXD05CgWthoXyh8jTjJp/DMH+EZXj1HCNu+X5Wf6lmincDcInvl9BS
Q9wpmYysp38H6l4kOMZXUEqTTdi1LrfXgUdy0L5w5CVu5JkRU3oiJGcM99E6Xbo0
5YyE7kQnxoydi1lCMcJBRj0LCy/k96/2mIvUQZjexCjuvGyH0pZ741ZZHdL4uoDM
/MM0o+bPC5BhMh4mIkiYSX+eUihORVVbOtifLNwtD0LJ5Q8451gMBG4r0RKXoYnw
uVS4tlMdrJmERVypCLRcYeoxd1y8JybFHF2oj/cVS4rONZM7260zlDhmUL6Mo8N2
FhTIwGKDLSX3WMoCh3qTP3GUWnnSWMLEcTksjqDtC5ryX7hrcajHT1TTik4Vr5lI
UVqYrtDc5RJTe8mMJ9eKx3mLPoJUc03jWMYGiO2i6ruuv7lX/7J7UWlrUvckLkoS
vPJYS39Do1NRNFwtovUcLblP0pHK+Hz7oInyPhzK3Iq2CKegaeb+wffGDYqdJtWQ
6ExK8MkFqi8Z2RPXmsg9ycHQ0OpPrY71ndAxb5KjahYT6JpNzJDuRT06aA+/gAZo
1jGwnnLKXXBYCDzyevSnR3auX2A53x2sghf6e3anyAICVtbsJihgvxPz+r1kYfCb
wH70oXBG76OapeIPwD4YWaE1SSv/Kj/lkejvAwp3d9WToCEuifUY49qpk5hoPe6K
NuwOz9qCvb0PK035o8f/kZx+g3jBhj2qDBChSqrdEF7x3u28mnbM5jmrWHwO6vdj
GoWz2dG0vS1vgluGs+G8XsMFyJe20XPZEh3bf8unIeaIyQqbarneQwwduQy/Ocap
Ader6BB9C/KCbpdeWRuc5zaWVF0Db1TSlyQXQA5sfdxYIz1hQwTnYhITv5S89GVa
q3X8jJ4WE1TbKA7AAoWDwOHXAMUz/imTf/aterUGMxki0ogNdRqjyfwCwpD9KsSD
sQq5MvItQjQjw6HuU9M0sXz2jpiCeZitsX1p4QZ9rH6RV0BeGT4PZ6+NYuRRW5+e
CIem4kgc7PR43UzHLSgoAMvQnKnGrngK5qkvc9IuyxJ8yAxK1bWJtp0QM7fcdmQH
X/F2i9USyNIwB9lhYdEFC7YZX/RvpTc+Y9iuJIezVClH74hHgeM5T36lyfGgn3Fn
Sr0BAsM16wLfXnKtROU14u5hQjjLLYSnpkrDbnyNNGWwPdtWfl3mclT88j4Q07by
ArFfPXSCKvis+Zx7wTFJ3Vmv7xdgB6MM3RULFNesyXayr2nuWcEG9+VBJmg4A+N6
13WhgRcXsa2wnWLe4KnByYX22PcehHoDGLZca+lMDOCcNUbxzcUNwJ/QNy0/rc/8
Gus/o02ltfhOCJP8ucJzzm5LVr1nNoaFc2OstAB1sWSs02eSDA6YMgrAmZvfs+5o
GDpnIRkH9hNV95K7jCTUVI4/cJQnx5trkRdefAWhAisZiShnESpye59LFBKwngfo
BWedSyttZ3XBd84HUIq9RnmMKxrJQcAHMMlIM0UH0zncShbdvlKkqvzdiPLNg8hY
h/Dai74B22l3z+DwhPrcBNhb+4t0/ZlYmpJOqL2q+8lZN076/N1IF7pxABa6rtr0
mtnf5z2F1xiRjMJmYkiFocUTDmnFgPdEeWO/Vyfyy4HsKpvRxe9+/wnF6983XjuW
JjKxd0iXvDL5Ij4l51fhFFrQe35fZJSjkAgY04sIPX+eVeIiilnKSJa+RCYZZZJn
oYJ8wPXvMroALaUNbTQwSKcihoy9BbGnAnh7jIIS0Kk+O3zULZ2gdwBADUi+9pWD
zKBTY0GREbUETKh8TGD7aP9naTkRweHml+dU6dmXImEtbML2XJ8BY9/fjtx6IL8x
DtIg7CsNq95jJggfl/9bq6XMlr6FnWR4CxBU6KpR3i34GsEwobIPUeQWpghDgLGN
xBEXYOAFurknKmNELqMJ6mFcIhC2qTWVmbmLs8RgeVGg+w5EasG/yIAZERncybU3
y9xiWVVyXhAroUeYa0e4RKUEnl5Ws5OB23rorcvjcT98u38gHZqlTH+ifSGzZK8y
0X1xB6ryTMMNxmqjFHKaPe/Fw3XaeSQdT9Sj9k4U5IF6W9xTzjKEeozCnAQQZbwG
fpyVwYEBIF4mU7hJtBIiNOq54wFk6+Q/Mqnuakv84aTx6WhXhns9qKKGDICjsNyS
Mr0qwY7LSGwlttHLSQHPpMR4klIEn0V7wv9PFf/rQBQXAEVHHbfo9OBBT6in7OhM
vOvYYuhOiNf1cRuonLgtqzlC88G9X5foCsfDv8sAagDF+/4KLYGm9oY/GrLnuuum
7BQFej167GTj4JF+C8cTcQp5YcQ7T6dS4NM3wo4cdKZblcuN8GhNwwcLjnaUrqka
oBS4ZiDaJdW0CrfiWwfWfS5V2tOZTH+QFR6IAdZ53h4/Vau61RJCBSmRUBQGUAxp
EMpqNg78e0PSR7+T+ntMg0UkAp2w9jydNCni5cSbXkPGgD339uHxmDNvYTqvv3p0
Km4HLgMP+7TNVZNv1wBpy+KpJFHiS1c1Ysp959lssz8ZJjMgt1VyNtxr/6TpfkFr
qlbkgLT/HreMGQJYmRq1+BQ6niSK1CDNZrzjFIxcELN3j6oe88DKeq9mMIDHAa80
bSVE++TRH45gLdbmipCixwBxwgfTm7yvQDQteyTDI202w3XqWa4kq1gQGeUq9uzl
udnwe40tzq4nH6CKkA5fQ3lUsxbo0NQ4seCq11rq+To7R+uk9K/TKt4n/OsVdmL0
M/ZFOHvHOJVqUKOu1QKAfp+7jgvZB11NK9QNoJDbnFXTbZxbR2dK24E0gUb1wMyO
ZCsF5jH14pilKrd+pQI5u9NCPk79SoJRllJbBbW7yuaPN9BtmKBTSNQobsjVmCto
4Kn4qondNJoDVYGnq8xa9IkCf1488xxzYt7zUrWM7H4GaBkNNQqqJpRhmKVfpU9k
lHV2mTQM7qy7W2cwefqxRlZLZ8BsXhOVNxnVGIknffZpJxibUQV+BnG7rmFD4eGz
mpwtSAPjhBMCpXleMFRj/yDcc+aIsTrhbGxHNrc8Mz4arRUxt9B53hyY4yn9Zd+c
u6wBLEMRVGiZIda8cTdbbTcfSV9kvDbE+RXzgc5sCZUWAeIL99TNC94H3BeQ0etu
xvNni0IOukSdrQ4ic5D7A3woWiW3n/d75dKw9WM11cvr+WNmK2uD1cppNBkyi7wN
/yQEKVK2vL1XigZaHKbykk+A6YsP8h7vbq0+wmZxhq2eushK8quPr3rqn7fcYMEE
lBynhYIqeQNYBRkLF1Q+7ioU020gRtKwogoieOZ5WaIst69VGtOMQBifkQbX2xJC
4eyY0udAn5usFsDwlxNU80Dlb23AbMOd05AJnQhF28ymZYgHr3yJjeWMZDeok54K
R+N3Fg3mhimXUBXwuPt/ZPz7UDlvwTXqPPM8YY6rDGollL1goY87m3KK2maMVIQK
6x5aDW7tiDOn5qOI4Fd38WclA4GBEAr45PDzLG1agV9Q9IjxUyWppGVB3a15xjUe
wIjG6MjMwJjyTMW25iJXZlwwNUhZYDXsEkWQPDdHd8qCAWoW6S/bq9zA45hnjkBR
4qlFggYPOhJyZYOJMgopBrY/bDL1MJnssmNe34eA5pVrWTeOsKIV6r/lqp+BH7Kk
8AouZKhR5grR517Fe5oNWvZEVrN59RsjyfAY3/JKKb/5OAhyj5jRzclzAe9Fw3xX
zNMxOjqJQK1njgNIYyF1IctvHZGulgAFaiojpM0shpZUNHqk1g+4CKZ+ACVJYLES
BTc1/hCXigwRR8ssbw4iI3MvfK4wdYwFVUabhLTPcdUKYgeet3AfChXVPDaj0zOg
hVQyldG14iuc3gIrvK1k0X824A0VjT/P/6PsiK2X9oMTJvoE7nDW6XELP1ZAPnwx
j42M2sAg/UPClgsMdqdIDogbwc1TfuKHNJs/0ly4gldJ+KrKy/fu/Dz7mEggeJ5M
mcFDkpLIsqfKFlhWnabIkD0iAXemEJEHBmT4q+djBV0VYZEr1+aKdcLyn5e6uJLO
i8xRV/pJGK5BDoDEnLzzj9X07PUcFj+r72BJqAgI5A+fHkPFfW42LAJBCo0VFsuX
L1Zhd5W8/QKLstSVKkYfjOIkqvsH6u6adtYtM6iduM1Omi2CMRYwFukB1hvkwW9z
l5WGBprLgsoOwZPgnc1QROxIStdGYn0IRKxOvOU5Ej4sDkG/JGgfIRWxeFbwNJx9
MDE7sDi5uOZIHhJbmbS9BoCMMLneMW+LCCDzFNR7xOCHp3Bo42NY8nFY8+GVaLTr
WKTgeu6c3x9eUSKLDfKd5dfgUq/ssG0CSpakA++LK2KV+i/xNurhEdsVNjbdcUQ0
2rVTybLkMaUZKDZIGvy828PE0u+DShe93pjF3Kvh0SCxKhiomRX6358Cf93SrgrF
qiTWKB5koaZXpT5dJHV1L1ynBnjQaVPpVZIGmur/AnTN/hSu/IEXHK2LUKL5SvpT
bktu4YGo68J/jpPLGdQsrx94gdHoi6ujqGtEZe/mQFtXMplwGp9/iKhYexAkoH88
5BZ7pU1i7Tr1AYl7/Uo5lhfs51oNAYotiZgtOI3bNtggc8NtpvyrpIKdEbpiT8lX
K6yZpZ+YL6EBfAkOyvtBtLmk6Q4J6NP5Tnm2Qk8VoJOwCiG8R6PN3IQ4qAtG/qCg
M9bJsyYTnE24+A4qUlvy+iOiLI7aY+nXzNQTnTL6RHXEV4pwELJehwRk1zMiK/ZP
3ibjrCzi577134SV2Do8gilPhsflDgx4SrNefnrfMdirhYbXnw+ZycMVxOFtkOPO
yPxKprbm4aYk2JmiArNExLcB4C3VVasBxmE/abB0jnFSs8iqDV9nlvtyTrvtOfmb
Js30LZvVnD6T9jqfsZ0U/mk0XSqVH2lMVz5JOKFDwyKviHoVvOM2k/NecTezucbL
ZzdzBR9PCYw1hpCSL/AP8z0cVOit59Ilpq08Bvn/0rj1jdOSmFKSW91JFxxfrwQc
YjyqMTU7SQXEmjy1iibvS41swtYu3G8fB2zGOvJ2YJrxS7kFYDyDFNMu6X8wfWu/
UOsf4T6WZmRiYZ71W2pJLl5yVmmJ8Oqci4dkN6JLYDEQuHNnK1g0JJz3jfJt0/gY
nQNUvSgJsZusrhm6TqTD8QO07GomlwEKsPjXiVdGEX857CRtcNeKZiJxTe9X/ao2
0jaC6FxrxE6GfE0r2PfIMGr+8tvbRyVuz0zXVqI4+HiEYQFlWUZYwJqgFY8fF1Gc
Agh5zJGDukr9v5CY+dFBAZRbI8pwPhj4rHI/WPcMtiSikkL/tRwygGyHCRTWcyIq
GZhzmPkiaSW/Js6v1f0ze/9j1rv6g4PsUhj1wJh72liX+rBIy7Tz6yGVvt7Ro5kG
czV91Uwz5oAvpKYeho17a5ot/G16FsHzKNs5kfGyZc4q7u0SaT5YEclYNP2d3ohS
edr4ROLBCBTYU+dkAGRHy9Azu8IEK/4y6mRhSzgqA06P8YnxoP/3z4mG8eSkQAgu
vieycAsB8r/b+FB10r6H4cR3x+HmTdALgVRG/vh6PrME04CpifS+wpDz+lyr8VoA
Q5+ZRCP4V3oERtHWatXposu7nBOvirwEI/owauLmLkorwk9VhQC11azl+nv8lW1M
nsm7J2yLaHGRrzI60quCReL6+mcQPg+pgFJprfybJdd11spoQNBxkLakZ9r48hWl
N2PI1PTB59hIOg9fSC9emvJdZ172cnK3uo6buCJ9r+mzOtM1uoYSSCa2HOUnpxcr
XzFXLeSeGXbqqXPtt50TJ4GWSksVu2kQ1y9FYduzl/mb7+pFB+WT2uKBOxzqklOc
1naC/yv3/0tEVB4GISqfXUdS/OTvrteoTd1HCxn64+LdlVjBTvQEhSB2jtd69gT1
hBw1lpGEcJTnHrUDatEaOO6OuddyR8EzJmyIi0+iXtftQKMNUBeu1iEg3CnB95wX
vD4MQnpIg9OJbjAxVSWNK2LoPdtLO1QEmybTIFFN4S3hiBE3lUIKTlYeVqFhfPgv
b2tx4Db2y5mkbSNms6OIBtq9ryTY2fHZjCh7pBiWRXxe1G/m/W77XifAtCOOBzLm
w+NCNkHiAvLMRw3FtJmGEUOeFocADeYfNtStbNocmkS3+bgxwLiu7Of/Fw1oPGVk
ICUU6vIYyuC12dgkqSi6jQJbVwmfDvtHVGz5HTdyhON2+2V0egisDb7LefBUPPgU
JAV4aNuR3T9XufHSUNmzxldihmyKuadk6bv8OgeYpMKAXrB9+ejkx92dHHyPsQ7M
Azj4QKwFMqWDQ0wPG6NEju+AdxB2jhuKmES6LL/LdjeJZLcL5GnOevHgdxD2tjhe
PXl5QOD68mNs5b8kYhdki03Rpu3YTVKxuT3H9hmpLjc17DYeq+O15KJ6p207uBij
srhkYDYNCwQ/8U+AeivWjTGXgPXLwCST4UFSe1Qoj72nXAqhXgM6k+Dht3hguF+b
61Dc9Wt8day5ClUtmwItvXwrOwtzkkT38EAlfSRaAEGqx6VhTLKlK8EvFnkCSMe8
WMxFhiWtASL7soRYxr52n3t6oRp7Jhf7GciBnvznOwRoCquMsRyrdVOwsBD3LXO1
GJ0uYK7ntCE3uGwLKRwcCJZKaBY1keiEocRurZAv8odQYF17QJJpeV0GaKS1X44l
rzG+BLPGr4oQdXw70djzeIFfp2JdDqdlHCVNom7rjMRswIK+LLenDj2QkD9HJNNo
5R8r13EctjCB99KoOt8HnBnYYoF6sXKkOoF6hjmz/WWOF57krSCb4a1l6mkQrOwC
psC5vRtR2ZaXXKvVB3aDp53FPAWgxaF3YvvJZv6yqEjOWeIT0MAIL6i0mVIhD656
5O10hilazps2zecnA3G4xhuPAM/g0jrXOSe2hMhauNdGUTHrSgsgDvXdcv0mx6Ok
oTN74ffkMhShskC66+95TZ+NqYB8MWIXS45iP1CLPfSy38gSH7dJ2goXe3wMR6yL
Bzr2aVZi3iYxOUhIAvB9dJ8uUvK0i+FyE0Pp5RaMMjYJl6bK4ufUfsPccQ+AwyBk
w+Pz1hZBkdUhu2ERishhrFWRegxfB9tNqme0rzaH2VTC8rYOnXZE+nidRk04x5Z7
hGam4giA/3NQz5Z6+4ewjuOxPHgz7s6A5OEIXGbmLSZSSWsFRyS+nLWUN4Sq2WnT
NDgV42tishcjj0/F1q+bgMsT3KwAo79O7gJTieEHB5eDcXYwP+L3V5nw6r63ACy4
qjf/zAzqP9ztFv+RzAFxsv71HADlhsym2CQPc9/bt368QaHFMpdqncW4kjJEhH3Z
XNfcbLMdqD2pIEM6GeD3WFn1qjUGtsNkF35FCCtWTJDH84a2f3NY4bqJVb0SJTkU
ciwvG3dlZbpC9BEKb8WLMQqjOFyb3xGUVM10SiWUa37raygsZ1VKLXNI/EdkOqeZ
zQpXnY0K9EeKgvqqlcpfg+Byuc+udZJ5r8ezXjRQnlQVxSOjSktMSgEMp0wWEwan
hvr+aRT/qfBi0a/RQu3CbKqGeVwjvrU0PlD2pSRMPexCyK7sfplcHkYXEpAjSzA4
hPQkuFegRtHO7Z/kES5t8xPZC0JcQmYO2vjVw7LtcvzHIMIXLBZydjrz3OcIvU5P
MvIQhGI2qvCTkp6+fjFfeWWcFi34Mbq3X9lX0yYD1VDre0VDMmZZDNyxwUKKNg9l
JRlOPNiO/ANqltMKptJV9MIL48rjB509SmCvAwc+MqB2ML1EHtrL9MZEvhhKEylt
CHcW4wJFVwl8M/teqJPJqB3tXgVwdvySwVSf1LX0UbP5Kaofb2WbyJqk0bKiJNuH
zjL3Tg6CWaqz4ODBqxu86zXjv/x0+wcz/z0lQY1xILeUXmZ4Z8B+GmOlTIqEeAF2
/a5OFbZNyOEa1pfHc76g05vfwsPiHw+C0mD95SMX57i0t4by61TwV5lWq2V3GUnG
QM5C2jdtyzTAup8Lz3NmgE33kmVs3tgj0XeAzsINnxfPaXpQA/Ey+K04qKRsZexK
wNE1qW9QpilnuYORp3hZaiLDSXzWqai09gUSvdFkqrct3kuPa6tH1dI48kHySQt4
lecbRTIb+20JO8BpWX/tu90W3R4+ZZ4+koS0m5ayfE1WAJUiO18h8i6sP/Eczyje
WgClaPmrAqqCy9eA2LAFzb2WzooaSlA+Vgp46/4zkEzDeAjN8V7gAfrKL5CyZT0x
LqQqjgNHufxgXSa1ps6156GoXqxwA40IulPxGH7JUFMYQCgcDI25VoInU5xM3/VK
QjheGVP0A5uG96igdg22o8UTif/cp7LmztNaprF8RsDC/0z/KpLl/ejI4sLd6hKM
6DRyVHwyE48rh9Sgyp4Ba4m7wxjAGbFEsqrL2ERf0tZjfnBKF19eiDygk7GNJ+bG
Zd8HTh1TaDXr0BO8+tEwPH+R99WgDdWmPHPZoe9oNg3ZOu0W4OzKKvXJDjUyQ4+i
OnuFcrx2iIOM1/4uE8bWBZYkStoHlZoHpe9pqjtcmlxw4z7OJXMGfG6NPFuyMCOV
J6cITYXX+cXV0cuMWiIpaFWajdqp1QO9k/YD0CTqJs4ucZn/OMeLiDcxJnFAmK75
e5UWDyVKGOfKy0uymniOUbppe5l3hC0mdO6voy/KhD3xqNKrwGZDlQByAMKHPzwH
Gn0MBG2Q4NzRnRcBQa2CbZaIaMz6M77n8Qu6uNl+rzi9U7tnqSz+OgE/x+DhIDXY
J2PZ3GtGB3mIekEP98ks0tI1iv44FV9vsYF5GRuZ1BTaDjJX4VqqRn3hGumA4BcC
Avh1JuFb7hsnIZLz10LZHqkUD3zDZbtQV41G+4BzLE1zSQmG9oTl1ypUprez3Upb
yrCv94aIpvfbh793iGYk9ZNMDs0iOOVGKO9LzPE1QSWGwNfxF1cDGyqsKTQPWfm2
z7PsKsEaAfR9ECNOdS1Mn78vAmKyMJKdROz2FJwz25d3xg8l+fMcmBXFcA0plOoR
EJdiDHYnNeq6JkIcm8EXWQ6mt58Jy+d0ESVkGKBCLmO6GBJUmBok0v4xW+XcBnaY
bub6FSOVGG+lfgsl/o8fIRbNyJqO01z9LsKQTp4IDdoN6RnMqJc8ouUsOxD5ZBKr
vOFzeEP3hJElNeUjuDqJQSQ5hQiKjcH6ITK9r41SvlDaPC9FM82ThhuSOd5aN93Y
p41k1vOkhVe7WiDw0a0JJHOk5zRAeazavpAWTrVqgRGSDpbRIrwRlLD4MUTP/Mgt
uGWmrBeTMhcff3oKXenEn7rJvNY8Oqoc+3WfBChxQ1bE+QKr2EFAoK99QcfMopAX
WrKPHf0ZQapQeX/r05K5EHxQU7jEzxhJ2NSEQNJy6LF7ffe+Qy6hnArV6ETR4L/d
VGLBH5JGc7wrtafh3Ny/0buzrxB89SHwh1nSR9MgkheFrelNvS3ZghKnIGk0IsX9
xrfN1PUyCNhpYuB5bcQU/6+FE/4aIKUoZ1q143gKoyZ0p8HVm4EFav/NDWCC+s/B
s8g4BnwRfuKIf4+KGrCgqbQzfFXgOMkwGGieBcCJfkL4aBaqLpVM+hW+zCwjUdfB
f/e4SPTxLWlSBonHYmWEy3AM/HO0Y7GWi5g2kNoP9CufGcZGAX/5XcxreN17hxUq
1Dl4Ztqb+8/zndOWY6v8FtmEs5cyQVGloRJealwoJGiQ3ju+5WtzREETlPnnvhiw
ml03C7w4NrH6vyLWtl5jBmNvYQ4qRK2nOMRjWU+QDEHtrJOgNaMH/2Ggmxxn8TsO
8eqry1U6r8oekg5yoKQme955zpwNN8nzyemWQkOGCECDpXN/9X9DDGSZtP2RCouX
XPreoBSg3uMLTNqn1AQnEGlgl+QuHl1+c61m7NZnUsoSv17I/qhBo/R83eEVp+s7
YxS2u8ca6B0vJQQVfbEmdFoqxt1WqP+CuF0kcox0Vrx1WLpsjp1aT/t099Nd2EeZ
yCe0msNQbpDHJ7xKrSUJCBo4sXkqMVWIVKQ3OewccHCgx+E/zXtDFLX4EuEGwWGX
SU69+oiU8pmeP1G77E8fmqTxXZhmVZ+7voU8qFVZgWFmzriCCcSMxU87maiiDMFo
G6eMzYyTU4GxlyYkGhMd46W2gwVYmtvHggzSdrBBtBg7tAvjZ2zjewjQhGDaCzv5
4oT77PCsV8j/QHuGUXVOgAm8Dt4KGBjihoLFVT8pK0OzamLlrGBMq6cBlaiHMA1a
aex6GSYYCPQb7GPXiMj2geNzcw/eH/WH4z/HSiHiQppjB+0RUvMHWWUt5QKZwA7+
BwfHLgiFn/OeLvvdp9MDmKbI+2RNrtL+YwbQVcQCKUOWxX+0eLxQNyo3Aq3r1u9h
W+IgK8rEJzhVkC7vX2BDDYvc9PjMpvAnbeXIWLFe23ad2k1gqE5YHSi+GSYI+haH
D7GAMwfG2yAJe3tXb6R5r16n16K3AncBPF8zqh4s9ZQ8vJd/Am2SZygycmqJjcc+
8NSkemjHwLYxRrCgbRZc61ri4Q4rgi8XMDIdDjHeBk+eksGDzP0YFtJDZyTY8CmL
mTkNYOg1Axasn2tZ4RnXYAzYqhaTmNVKotqtCAQU8e2c6HvQoUJ8YcULxHxbrxez
1soPyFFf7zIeixrkpthJBykowGD/0VDvJjIbh7BKl5g7wJUFdt0eV1Vq2um8Prwd
hJnTlD0f/1YaWYUcnfanhI6tHdMpavZKeHSeJegWvxyTe3q1y2C7BRi3/N5Pk66U
Fk++sQrQQEJ5GuT4p8te+LByvPyQGYRdVGsjyH8x5S8486Bvm0GD9QKdwMBqLn7+
5eube8oLTI6dYxcxCaFeIVv4elMzuNNKgs88NkdFIWNK4DaeSWrYE9ai9QI/3CfU
xMyuQNkndZ0hntHQyn8Ct6s42TbIghMKE+FlJty36ZWuXpzJklNY6twZbC40Gbxo
xZgGv5pLoQOlgSQ61m0qCY6zLTtrG2/cv3/YUzthYtf70iL8kXqrn3m5nG2H0dhn
2u/LJSdwcscdh1KIg6PIduqDsKcpr/IvUPJeWBlAhUzgXLiBSBBWbgscAZ0UuORk
MeQcpIKL7xrPAl7lmJDKy5Ldnoz5NtXZAAt8J4xdwRS6sUsSS+CA6QAFfwlEdvQb
9VMHY0cOqNKBu6BzmQN2/AAl+u1KOmJyvsIXMUrgiVPdqs6ff7gGwcV1nLqWGvHV
0MikxsteCGYlibxSnFyBfHQmvzsZx3pQGryx5rT9HaMRKN8S90OeQqkP6orVTVUk
7giwCkQhWjYVm6UuLeesh1rMAV445Mm99zzjnckA+7vYwlhetlk6pgJ46nxlpuVh
uO8phd8orzDfgg9rPddRl1eOshLxQvvK9qYstrRRbM2HYwrJWcSWNEVSQz5S5ztr
YMsaS6HNIRHpBQtDwpsENB7U69+NiJKtcmfSCoHIeB0h7UAjdPll3NXeSQ3kLEwP
E5v7tvZQKBZ4vmkBNNlQYmE2kwsJXsBRrA5gGxWm0ue02kHda0XpheLxbwxNEzKu
ofs+UPqr4iPTCYfh+Lty5cypufUHqRfxgQZdO9ts9+SFQVab8gdLk2dvDcEPo5dG
5lFGkbo1ZERqZ0Hk0EJt/NCxSD027Lsi2knIdW4Q6D6SCSpvRPctNnF5966paijn
LyxTkJENAD2iZmVG+JLnXSIKoHWc/4rqWuhn7o605tz9pl1NagXe+M5qcSRmXfRr
6Ow+QBd6b7ew+WE+lncVkO2jL1xnZXWqelBvgW9btk8fSD7I0HX98MRbtGcv7wYb
2f//KQyFb+vHSHt8GZ+nnVyZdOgj+5zdLbc6fw13Dz/g8BQ/ciURkLaZY+2JMq/j
3ZCqsYAC8ZHJvItzpYf21yLH7y7ZJN54Ge8xP4/le2l16GT7lcDx+5s98zemaBvf
XV2dRVrtzDpmtkWHVGpXD2eE4VRQlaLcMYvzTUBDNkn0Cbhwv4ensUfuGPE9GmTw
82RM794HBK3rKUiXkUOYgKjyMXWSF2hIlM1t2MiZpOxsqEgrmcgf5m8cRFPaYPYZ
pRpYY1zBqRRHMBCjxwmRkhgS+eEv5WA4dLUmhXub4OXCCiju+dW6wK4FysWlHtO6
mhiciEpDxRdBnD+FEChx2wfR3BZo2TOQlfoUk5hw/FIQvfwakV5LDU7TDQbeuMNe
9L4fQSku6efkj6W6HrD9IKab6UqEElD5yp6PDrXmCLWqcN5lwCD6lrn9I+NznUvv
AxUSEDY/Znw3MhPZ/4abrTCll3J2RnJ1+6Hn4a6wijcWyfQ6Mqn+FLQPGdw9JMZg
2Ip7OyNFqQi9Lt+Cw1AVE4i4K0R9ccDVMMWOUO6b8tGqFOXg1L2dXvDzt2n9HD3M
S6A4Ed2NgFIAFhsGNDZ9rM1IgMFp5hZpQJd5FK8Lx9cxeDJREZ1UJl4ENZnJB3Mk
2NxRyUvgc7Lb6wfTxY+zX30Da3ZgRpwddDc3e5b9tmaiUIux5gwX56Mc+i9DB0n/
GvLp8LJvhpBcbewjd+fJ7J/eRxBNdS/6Gm5t0p/d0BFQVj9M5OmhGo34Z7juboU1
iaD8Z2uD6X94wpndkbhSOcbjNwWMn/KghSZDfGNcTFK5zjGe64CxQy+RYFBefboP
I7XTYNHE7RRXl2mMxr1+H1Maryi9vKyPtQx5tm7HMo2ubscSGLe413oC0Q25BXjd
zw5j76Dd/BBX7AnCuPnwm2NVsJq/7+0hvncxs2QajuiTSFZczMX2Jl44Vdht8ShE
XdGz3Y6Mzyp8P82w5fsyp5dwXAFYpo8+3QTDUn3dp47AkpMUHilcLQKH67nIwQlC
/ee+ITktVaRkNRhXD2Ngv7sl+dlQvQFWSXFiQ9MSUROd7uK1LZ7MZZLntB35+5pl
D9zA1XlVyqTtB9ipC0qsgJaZ5xUMGmgm8yFlAezBQCFjy6nq2YQnZQ8YlgNRqdIN
NGVcoyWMaKJk/rkQ9GfoOgsFCcYeVbNRAWZTxZ1By/SPmJrnEeBhAUraYARHOM2U
XrGpw5KJOmU7T8Uq+sUn8CS8GmaVdbS2mpD9aEkogIXsx5ph9uUdgT7x9UqqOZB0
1I2RKwp0PgIW62H4drhKOCqdz1w0Tmb9c3xUPEkEz98HwdqeQJdb03sVsNLbX3xq
fDKaoyY+aSZo1s3m8f/QDGD4lX+CE9+qzs9gGXax1k6BBv+von34anWvgoJa1h/H
6tofd+vTtTl1WdWAqipWAEtcGMNFQGrVglocQleqlPOY1fUZQlLOsQ8AcSNl9Pjb
9rbdIc1YYbodDN3bnUfrqZ3i3jX2LdYHJnDWaKgQysKJRS7f2OaMyCD2dGs3lHCL
S+VgpbqkHACCKetoRbT8Kk2TpJyP+5orHTQdVB7o51NLZ4pBgiKViOgbWWAQ0e9Q
+sZd1TnLFlcRNFSYW3W9hXHtRn4zaMX1voZSUgl5QzZoMEh7uoH83aStQUBIAvak
9woDt49wedoN3FtqRp6RimWkfA8/YvvNxsARZi5wMIVz5zTvDtuqyoXIFfSvd5A+
wlb/dg78lFQygIOT/4WpDgYPlcEZC3+Jgj/gvMiEu/3XpK/PVdOGt9GtoLOXIgct
HOHQlignVJnI8BOjy/k9O73i0uaDenTw2PqHFmcpCSe5X5E9O4Unyv4kpBdS1X/Z
QJ/xoS5024GmQha7o8LxQ0X5Cu33iH8n2O9eZpXDTY3pq5CaxEylKAOf4NdRggRH
aLXUvKFHevN7tV/OByHaLj5x6waeQGtitKSBPL/l4oWQg3bYceM4H1qLiFi2OSgU
4i4cdhiQs2PzYJS9cTghz9FFlxTLft6xM3pn+x1ygTXFGtigLB7FOFKPlAYKfBu9
DIOjY4JhYCI/q8CFuGVhUVQlC09DXeT5vrGbCGU9PUvxlqsfuQ3cSEZLj/iJCgHg
OdGayQUz4gvF/Lzkf5dubNs8l9E96rXQdnMkuycr4oB9OWFhonYNO/DzWZJcmXgS
HWf5kGskqR0hoSYYhw7DrXwrPFKEugOe7PpdeGr1h83QWx2yDM1cBCPClfMtzZie
LKLlbd6oRU3S3XofRvi3x9DficIVKmDD/8I3/rgXYg4Y37+sldGALA/nE96vFXui
+9d11YVBIJJTOTDCH9/9i/qjmuTVeqnSdBSh5vT04XNvK0TjpXScCCp5p2VA/xhA
O9WETs4yDzSs3fW1JLZF2KR6KuobSFyo6nyGZSekCXrraNeO9xnwWQ//q7RnEHhL
GKGm3YZ08xtE3M1h9ugKLAMtGABCvjBAJe58ttapKsYjgNzLpS5BuagtKWPR3ume
uXo+e1nDHeK5glVcU7Lo8ikkKfA+LByUI/wSRjmKO0JX5lWVVpmE1Jj623KaDEnC
mWJZbXpRUO9eaH3osOpoq46Fn7hZ7X3BYuTKBJjuz48cFkf2+rM0wtr05F+vhp5+
IlcrnsRXMLvOCwOwoemfyDI2gV7Rfxm8U5NAIMeZ09FNq+8rdppNUC10VqVwyKMh
83hEzyMy3hseuW2C71beBdP/CUAn3hycoq+zOIt69FA/hld2/AFt7AzYwc/IkKWB
pt6LFuK8cJH3S3sKtlu2GA6FuArEmCgduNHBKiwxTTUJ0b5BLQ8qt88zwBuvqz3G
oCxK1Hbo2GaZ2yFRcPH4mhgck2fJJuuguWWOk1K6fcVRlZxucAVblHOMBXDwHvYA
N5upeDX0Tbv7S7ng+STIRQ4mz1apzIOQESAUrSQbRCr8o3FptvEtnye4cVk+xWxy
qKjpgIV2APc7ctbOuROSyR6OjMr6d6T70Pcg+sAgg+pZQA5Bwy8yl66pUR7axL3b
fXXct5Qc+1L7qRXcP0Y14BtSuBoBSKMtvAMhbxtR7RP7B/76mopzKX4M8Q1ZkdT5
DIOL9ikbyp9n/TDZvS8lvWAPRQwI4mZTw99y1LmDDinwPJWe9PwNyVPfdTqACgfK
8yUgme3kbSvW7EDKA1y7g1+NZXEIIyN1fMcwbYQtVqZlrbiJXeZ7IdD0LEhiyhr7
/df5zatIVJFosjk4o66+Jtckuk5LLIXudDfqUH/DAIZOR+XkgczTCM5CFiv0lTXH
ZbRqxDgu1J/lsicMzl97XL6Kz6LSejb4CxSJJwFbGUTHY64x1p+o0hxdSx49k3yy
8K+feWZ7+Ax0Fk3YOYMgZWp4r91P+j0SC+6AsO6RsT8QZsNXF/dSz9Oq6TL/hrL4
OmmDn2rbUD47ryyd4NbcGF5Y1tu8uMzC9Fxz+h8jsHEDNDZ7QFzqT0xpqBKDl5wg
EsMbld0AoSldYf6t/z7KMqzzFMeY8URGl6KDhEtyvUAHmraIA9vTrcaefEKaf5Bs
40BxgRBvfN/ohCNcG4n1LVFwh0dOE+I1lXvqrQq39LTCBgmVawUjM9o8lLly14/d
+oiWiW1gpVVdgELxEIrFW22hfIpxaj3W1f2Cdpmibw+RsZCu5KfguOdNh1V9H/y5
a3hKrOlJdwBnMKF0RdbMstzpKbwPC8aBp7lBAzW89OppBOGn7F+JVkilzhBvBKRe
nc0q6/q8CgqFuWjRzmPzBEd+l9I1bvaCic09CEFqnEZB/YBFphiLjRi0mOgP9Zw1
Wvtl8tsafa6iOwmnOR3ytOdWuLugS5D+o3Gdb7M1HxKGQjSLLLCJA1RBYr+t/ar1
8p6FFMA1L7tkgYd03IqCvoTMuo4p1yCTUz0g6Ho1MP28w1NzGK+SKytlQaX3tmdV
xLdmJmU4qIBzKEV2KJ3hKCyJUS6T/o+yR93kMGXFhXjL92ftSUYRQ0mtX+d3R1/j
bUocfX8YUGGjSAcKR7fzXG3jHaKA9/trHu1CJLC2OkQuufglv/SdJ1ifZhFbI6/S
7howu5RQa8+G6D7RsG9sm2tH6mYQ08Al5XZVufcjJbRj7e7A3Hy1EFXDqWRVr5Wm
IXDtltD5aodAXxCsuh7cEJG4LZodRljLzgWqCrn9IirsTLlZNEGqBJz9ZZUbi9j2
WIwU2NkoBr502N2+GQQ+oi5cK0vY0bfcI3mm/z2tPMdZK2ANNbzY7GoNNmYUpgd0
DVU5qUZUbm7mDxIGdv9YzaAXNmLB3J8TH92oMgQmnF9TLaXlZ/L7wzN7qTavTygn
JEN7ODnQ+mmYFIAFORcwrBQW9ngqz/CXK22+ZbHRJXmsp5JjsS4tW6FDpsJbi3sQ
g86hmAUqAoPK80RR7a6QU1r4aFM77pZq4MOSbNijZ3A/rceLr/V5Co2QhxAMrVya
IOiPuVA0J1WBieBxlF4pmLTyZDJ/5jqg3HDs5HN35CJto23lHoFNwZputgZMrbwi
9NzLk3OlKhbGr8BpFbrnxgeyQoH52wuPwHyuJALxdq2UahgYMbNHHFlgAGA1J9mV
QJMRHL7W9R3+okJgEiXL1V9TnNfoA52flTP8RsQF0rXVM/bdiJjxhgt+VDhErs9Y
wu3jx0ZjeCpcy+Ov/YzW5O2YunIREeMU01PZifbrI/glC9gaRZnOyN1mUt3Pg5LU
/gKX5d1ZQNUsSEAPwjBXIIaJEhPkkda3FKkFW2Yev/fDHOF5mlXDD65ZA/qh9f8H
658LtmjM2SZsuqcE3lZ5In0+Hm+Yk0Al4GuR/PHRV3LTYII5CRxFXdWLYRjHo3ib
cjbd+pVzolcSr//jo0MisNJqPWKs8iGO1b2Ou+lXeFe4zHjfW0cY0BUCvpTanbPX
L/hH2rd3JXHDKl0XfJOehY1YevEDQQNyR9LlhMylJOnaFyNFCacpVuSi0yqrodBb
T3sdWFxNe6TLFOTHErQxH4g2c5N+724z0jr4TyRLzK4f/VexqxA5ZCYq21opSpqa
P3+2D3uUjXogcsXBGH1ieun9QwcPjXH1t0lT/WHOdjwAH89XO0+ideRLLxmLP8RG
qy/9p7AQTE/4ybWuxPOONcyECnxT2FjijiekUEvhsT8gN3T1WlH0Y+A+GaUx0vWO
nwT+t/gXkqGLkDw8szeQPWtxEvvNjqG/UtjQV7nQAhAlu8XZtHdto8kqmNayigSw
Xphj135A5j+z865JF5cpXaedHPg9gCecWHDqBcN+rR4a0iLtrLWBiguwkDMSaJqY
v5g81piUgGhn+TyWiHiY3OVdwzaC4zAc/iwBKd9uD2Zg3/L0EeX/IU3FnvnVlwf/
czXpKhCGbopr94tQ0DGywRSZgKFFNuW7t1gu4q/GpVSLEE5wqPoFxp+3JRfYCXbh
2gjge57YKx8cpvJ9Fvam7c9JIoE8VyM/GCXe9T1BbsF7qF4EyLQu9jCdPns4Rs7n
LLPccDvWigybrUsmk2XFfa2JnfSq+guL5twgxUy5c45kYFOnb5F8h4yqZsUg9Jbg
QSkh8rpkGETkN469mpMGH8BmrAekBgQd2oxabUx8FDlkuSIO2rnccij6zdkbVoTt
NgkLid0i4cwiYKoRPrWPDa8wIIvr1brG5eMr9nJ6gyqBgHFR2po3Xz93NPx8JfOT
ImclVYGOPJazrwrL2dLB28gLcpP7YgJ9Z/Ri1qWbQQSm/CjCqFRpoLpdPTexGR9v
GhtG8ujSKlx4TgeOSWaSbQsKbnm0Wv8L3HHDxjyUlTJaR04HqhaOHf0mty8etlXP
F2doZJu6tSOuXRmj56Ceo7BQylZLdZUUiaRvbNc/wdvjYaFeJq12/AyYkAHYegh8
rEX7m6DW5hoCEhZhnDJMnajcJrLZR1ntSK77Pm20JRqTMM+vAHZEzxCrF/YsaKUP
uCRbWqP5YNDe78FXcMOh92qyVAkHrDyWB157c4kmVn/2YOqjM6qrU237sLKPTVDn
lJOSkZw7qkL1cSmovRW+YM1SFb3atNSut59XuzHJeREduVM7eWGsQMcT0rsaiMrt
xzT8Qh6jpK4ARTPlHYt9XrdxbNs0mEXc2MP202gw8TJ33kBfN3lYNh3YkknCoP/w
N3ZEVTRrwzVbfn/xdObAT/IcSVbXTc8lGgNV75F29ZwVYKSRbtTK8FY20BvzAwTg
U9iyBS/8WcqnwRdEirTq/wttyjum8n5tcOzJK5cIjDDOTEL0aTinL2D/ElZMEdja
0VLw9S1Gkg4PT/0SgstCr8rkV/UIpfeKnqhH8rIDVUWqzMf4b0ydq/ZcwDUxdAai
VlseDo6j8xurWVLugaR3qfNAErM5LjYwVMl9sG96RiJusaq/c8072seDNg/JuJ7+
mffGzM2yfRv36+4CxrEpRtJIEZPn5ONdqE3xQV0L6SZwa8Nqe8wq7AkwEAeSODbA
hN8VkYjWSk3wF0SHjSPQ9c0tNTOgnpRUBUVF54b1EIa1hhSBnguUWCvIOD/EFFSz
c+a9FnGRN2xgvPr1klG3sRj1OvBvGVQvYjIvnA8xxKUefln/s+Pt6T8NtyWyUzdr
ivcUfANELV2bgM2py7IBRoHeH1UK10lEv6z2QqLIRfMf+oDlym43nYFSJ79kFf98
YVPWPGUnU7R+Ks6GLiBNQq2Q8PLJSDYWf6A9utfqXcMERJYYgmohIQs0dlkJnkEQ
efxbYG8LZicK3Ruu5fde5Nb2b9PwuGrDW+kSci+UZ/NGfOAKoM0LjZ2y2YtC2AJO
QwkUlX+t84zE40SBOaNot7+tMizp4okjtQrZHFbfz8NN3L9pQF6xxZwY9+s+r5dp
CAMwfMfr+575BBOddiaZUPHv284LvSYXzwNJV4iwuF7k07Y7QXF5fKgLudKFRGn7
kg9foeRVBtNDiJqXlpBKBHd+bsr5l66/awLtZRAtSQuOSr6exqh/gMfaVhDQCnS2
2ouF5lXQ6ykzxo1M5as/2EmMCDdKD+dVXcGaFNNoonWHGENPi13nosTp9yiAOVy7
uEvkiWR8gAG8cA2ZPqUtzC3gN70K1s/5DXAcNrUGSyK5aUd5IendsX3a6Exwxby5
RC82pI7PVLf+P3FgWpk5fAK5P1nQG0hy0lz7Wif9FDhNHqQ/BH2kNywl4Z/dVVFj
sxOiNe5NBgdzLuR8onXx7njCdHFsXUTDnGQEUz8jW8L/g4VzPazWuIwgNDNJLf0h
iGYbZB/RrfVpJAtj5jb7DW1Sd9l93PXZYGLxNbzpcGNCnfyN1d/UknzHTV3nIyj2
LX2dpQ1YuLiictdN6fGZbU2ypU+A5KJAuABrDgezl6WuQeICf41GtTDMIeamUsT4
7KpXmIroBi9yx0ikJz2fyCyJHa8RPeF7XiU3680RBCU3qxNtlpzKWZQsq3n2mB1v
hveJm/y9BOSC7LnXOpHAW0yQxz+7NRkrz6WaSHy/DNG1L16mlTeEf1CNnVzARnVf
UgLKzK9q1bYHfRV6bcDmHlsgliZk16UmZvPe3LUhGPONQJCOHCujuvt375h5PxB9
7rAATcjC8FOHgbfGO3D4VkeqWN7oDOprS1PU3CDYaNKAtlC+YES0/Ht33l+8e3c8
r8wtvS0XiWk1SDPg5mOQbI/ETfRlocohm3/wZADz6FLwhrheLclFYlK4G4sKM2fo
QIW/k0/afeJ/cdbc1C40RcuLNotgtnrGbxrJE8ccYLuL2RClftnwdYSKipXef5/T
iwgHecht4cXUVJe8ngX30BziPtph+EGvWPipwraL6ZymWVtiGXEuve78wiYItdjs
30oxP69Okslw4s6cUiPEvK8gS9JzJ1EbDL7MwhUehTV0VLZUJqwms2Ff36R7fPkV
QtM8OcHvxHb5ZhKsIYC8XK3JIIMB0oIgt653RSz88WUTxSf4EECra9LoVin0+dDO
QEjAc+G2RF2BvOBv76YeoUs1oKNgS2tufVRuCGPP20VW2NlhAAxey2JU9r8jm38/
7vELorGuPQbW60j+oBV0dClxbZvi3DOinWTO+HYU3FhX9vaDp4WKhIGCzBcSd6z+
mfbNnTNvyCLx/uGJvynfRbCUw+QVzCxRVWaZ412m7M4upheIf6VTKV8PiapPV/LQ
TuSkNOXXY2mug8AaeM9AOvAEKJiYHTp3UhYrrgWE8DAHiPBnJnBHK4xGTjqN/zwA
fmwjPV8uhmcuz+Plv+ck6wYMqgq3TKEEP26zDHAX0qP9F0B9UvGsLjg76LFEkUHV
cLkadMWcyLH8dt15X8um2dOw18DGy8bSIIlqdXS9gpAQqvgH4OuUYf+zTiI5EKyg
UWjXNJvxnl3zfJH7svyldlzWaaeRD0I8tEIvSUAjdHMYjLDMELAJWrPLEj1PayLl
dR5SZzFnHWWjsxOlwefy5ugmOVadpuDP43vn7qAm0cA63kU0BWVjw2yGb8+cDnCn
m6dqbE6L61KzKouG5zDlZswJlbYvNSgNwJR9YzISQpsXLTl3OOeCm6sgXFTZblDv
uCajTtvW1aWdW2Bw8Kgn4T1X1hvMKAirlO3EbovEPTT1XRWllDosDWhoWdNDi6L2
yRz6aZoMtUBeFKWAaEbTM51TismM/EjqXWsKgW60Lr1H0nBalDxyEjP8JOwkF2By
y6doaH9BH0Np16IxXiEFT6VlEiHMGP11YaM7sIEb8G68dyJ3CB83lZnUQ2CQ5+Fd
6xpwT5mE9AFDpjQDMDkJ2L/iypROVAF4rSJ3CCbgHF2movM1/Q9PzUVYoZS1MNsr
/K4nV41KQPQCH9V+lRGBD/pacEAxgW/3fKwVVvK1uxEwrVg/n6J6YUwiQOiu9sXx
ddXFMGONNEvczT7TjLW2qylOY5J9jLfwGRe+FwjK0YzD7Z4F+hnG+g/DDVVlpS7n
ou0RP+8YbmAV2sW6gdxYokA5H2pDJaC5432I6ho/1EpaJDz5cDzWguYgqruANJNf
Yb2Ux6f+EHZpkLwMl7uUnjPvA0j7fGAgVrZSeYuzVMR/qQTpmvYI0ZV+WWuYHz3l
pLUklBVHsnyNfmeZ0GHvdS6kAfOgTuSFSeSh9++k5hiKXZG2XLOsH3uDpMGSxDF+
bJ2Jk5pFUds/KYdih9FN20y4SPLtBSOoQ3VLax9zlnfIJUypSpR+qWYOPgFbmv0f
lSGdiQw2lBMmfOp8T4tN6WjeRLq6XJ6kArWejdnQ0HIR3v4sdPD4Na3jmjCEhr1i
B6b91cx5neK9xDhYxJ26KnH7qOe/OH8R3aEt21HOkzXgUaO3B6RM35aTAWnZc01T
ITDlyN+IS+w+pLyV6nf+ubXXE37nhu7FLAT0q2zOjMyqCA25vCy6y22KD/anlwuj
ib6KQrVmILZ23DVk67wajUgRbDIdvLk1D5Rszz2Rb0bqYSnNyKZgSJYf613hTcdX
WwiUMOPImOTXxrBbQ5WuJ9LNgwTc252YwLj2ZlpRZ45Ayfz7iQoRlUdx7Eat9j4C
aWQNQSrJS+RqFeWska0p0hFmSnmQmficfN+r0oBy+6e1L8OYYoKoSg6RICRwbSps
xrYFF2MvgF34MBo5hEBKHi14vM4zzo8TDhmKmZLz0ZDcuVMigdjn6o1kaL6GVjaf
tNBqLwbcSniuZkOEgbcknYCuJouFlJTvOM/OKGcJTOlr7ed67m1l8XhNwe/OZulH
GKThDN1Ne6MMwhWqFSZ3ZYraiCw16bZ6NfuJMuDJPTGnySgledU9sbrs/sDComtD
V4oRhWhU0OyhCF2adjVh5+QMScmN1FqO+1x814Jec7GNGP8s3sMmxbFwTKJo89tJ
MIfHkdy3fIvAxiTHZFHAlWuHB3XUyeuw45izUhWbJonZnmhoSm6qjVOw9z08VCAq
R5IjRxn+XQCD3CXVbOMQ60WNcg+oVEhMcLwT7p8WuTAEQJvuJOpLqKrcY3/2RcPt
70hkyqCwPF1xp6jGVIWMGrI8s6zHGRMzgFv+omVCYSO+EEOBt4KbzZWTZIXNQ01q
YSDpZd6EgKFiGqJQtEetZdxT+58ABxFizIoU5ASR0vUPyganSpIcxw2GUTHd/TSz
NDhMIkpibJi8LXNO4gn4yFpMQf4vLAeazB4n7lf0JGX9FbVT5SXsmgNQLBPy7D/V
5uvni7qjAJgenyRWX3I5b/tmpFHkpg/ewawS/kezn/BEo1cn5ODAxrqH1OjJvxj7
NW3QUXTqrirfszoiBTi2eKvOhDJFpDsF6bXyQw9fegy1a5PYci4PpXXuktpgXx4c
p/oP0w7Qw0C6kP//1b94FOKHddgRqPkejdDsyt6EJDaSA8R1l/qCrtGuFySX0W6/
Lgcwe/+D+z9qZ+aQKfs/1YMepvL3Nsv7356vgvDiTQ6L+kkgkUoDUpPE9kG+mOxq
94w08aaGFcyQGbrmMSNf+ge6MDutkd6FvyrSMIoyba4YCj6RJzvlgFDg8rab1fa5
IALBWrnkcbgCTh3envVjdKQ7AmsW0NgSEkC/mb23q216ARbEgv0vNjv3JfH8FD0G
Fy56yxcPfgxAHgzP2suSUQJFlpTmcc9BLUXELO/ifwszXn7hsOI18kNsetQAvUBg
m6iylGem85F4RFjX9yclfTfgOJNjKxBwC3MqN0luaVPGcBvKrAYeMPeRle/AHUPR
C/xNiK7kutFcUWZYeXEy69Mn/oNbFnOtTiMXiQGpKz/7aqN3g0q1yZsCF+xkqBxB
UnAnRYZXTwDjVtiSQvrynERxAru0L00YGvWhQ6TEa++hnr9A6x5Owwfh5Q/ZiLKl
V5+8nof7+xKehBRzOOmmcFKW/XnIpF4D+TN6W38LflfLuakV7eKy3szLHw8+LcmF
LgSzcYxETDw8W9vG+HZUFMQ6hJl+RGEaXlT3K5HqUBK//WnzAHFtFcyrDdWExAcM
95qDqHbiR8mEnukdNraNF/k0p5mVZOYwOv+fhUHHPg8cAufZDxymWyLB82YHTAnd
L8ysfdi31i0MUs8jWwlpuUl04dlobhfdQGAJJ+PFRf7g7Gx8wmROqsTEknljpLR/
6nbeQUyAYO+XczlbIcL6FKGu87rjvPmDWoF0FOM3KLx2+3MbTTmUuxKJD1GgoceI
jlsBP+iVT38fjAUHmicXv/fvKtP+dt1Qr5pWB0oSW+E7xY+gXcOXLFQNJNUGeiFQ
RiA0UL7gNmrv25aCQEp3QZ9ZLD7JkJKWcA+O+MV1x3dT7bZBvxuvKWOhfmUn2JIS
W1sqtzCcYsv1dITH6iEFGWiIo3CPwZk+StDW3/XnIgKvfNxgbY9ZKQZcicrnjgUg
fj+dqi/NSU3mDb9l+BXtbwT7Em+tQHbTDLhFneSdxUB4+SnNy/WVP+k0ymqG95Eh
0xiYvdhH5wdBXrksa9BmEjUsSDcykDpNOpBntKKnuexv6zlEEZHpJRwqeBlJ36Jc
WFTgSq23wF/6abCM+iiqRh3vq+jDm8YFsai82IWmwCGue9dL3AYSLKZ7QS3MLG5s
NImBnxdc59S2nPZDpCBxZiyevlWM5aQboTDZ3vRlJScuvLA2KXJHqQ5QDAN4I4GA
fdyBdAs6vWhP1s9J1GsRqLNwsoBPnV7SbE5J46vlnRF4ZI+T0XuvIQvKQOYQeE0B
YhE8IWc5ZBI71KJEyfhErXCptEzE5JRlGMG3XHb0TMTdjjtnzw6Kux19r4Aqwj6J
aSohQ4zpfBJy02iiFl4m9952mb/ZO+uNyqrW4poR3M6IA7efG37JSmicQ9DM+klf
PqFuI1f0z1b5zLYTf4NQ5GW0mYf1TYP25S1fsqzzbaT3c5CQIqBKW5Y7NlYgSU5c
bMg3MPMPykGrfPV46VBH2AgIV4tLoN1wZWQAdR4dFu941sOSyUhCCQRcM+ZSOE8Z
WTV8CBt2yiOFtrD2kmbsm7Q2KYhx8ho/jEgcejvVB4xbpn6RIl/vT1BjCwou7UWp
ORAFied0ZEH2ll23x8fO89HAEUPq7mirktxZ4hvowXQrMnljLnqwVh4XVT4SeFDa
sOaLXc/4oWbJALo8uOPmTbcTENOO6XTG+NyTSNeE1wqno1CeNeoEoQ1b8SMAFNIE
qPPmpT0OCmZU7r5Mwv9RPz6ohsnXShhqluI6gZ+Pf7xphCgkM5RePvyL61ajwQrs
FYA2oq2LRbezIYweLYvxGbk/OJCVcX/KYp7zuYJPke0vk0BUOnJAmjELUolSiZw/
HlMJI3dSar4lUyMqn+WKxdb7/5W+PZ3SeBR0JB4pm7/wMGUXHcr6e46tsCzmL7UA
8RFFOCIjxWMNQtQDIbj6tJsfRluhPZcsje2l3Ju7BWqfu1ldQfY96Mjkpswloa/s
oPTNuo6NDE6tT8YZ2A8AhA3szgW2gvIhYG1k1zFWejD8kJTNsBY+DZnRJYBQm8W8
zSnKKn+6Go7PxWRZv5KLPOQvcM7hrJDrAhc29MMFMFtqaDZuKSvn3aTW5ftp22O8
kZeQo5+YXVwjJdIzu4xv/NfVpQfcLNORtIgE+/N98Nbhb7egyKbVbG9vgwPo4F2E
soYTA8qko1HB8AcYO7P/srd+49vcJgocCnWrg60/xK7PmH4F0Kzsy6MjYRoj4MES
rXSHyqQ6y+KmWZWzTVqZV+B1iA5LPSRsUpzeQzqIiAQERhqbG00PhSnoqUWEoghN
PyM2JBDD3na8r9Q+fZFN47JftZCl8VoLXS27+ycS2PVmWWlmiBtcFO9iFRDb1zlH
9/fFhXwygoZSpaJKOn5Hhma96mlrByDAlOcpi/ylDqv9YndlK5ouDcqUuIuqh6yg
1hyS51A422iHQgFx87sKMvKUMn4vyZ6qPm6tbJxZfzKPdotBMJ4hl9MKGSUFtqEI
USryWY1sQsX3NDbCEjZv7AJpvIRWj4TGNEwUHQE7OZly04sEqzfQvGjT2AEsWLpI
ZSQidtxPUG73bYQ5xWp2XQ9iudyYt3/auLMhapLpNpvwLFqpXKcGTsqAbiaqRpJa
vlY0EiDvIFlKGCirPL4cWQft95MlNAteXqj6PY2hGaRY7MNqWgjccnJ9tN7OgejD
D93UzLJFJZYW0kJaflFZTChO24NEgcZvtRUQjp6qK5Rv6APm5cUSKvVz1e9ymbsx
kb+pYN/Z5absnseYy73nF779fz2A7+moVNk+Y8Ccdp4t1nt5jZL2rNF4eieR0nuj
OvM9DIjf+1WkOATM2tM7PqhCDzozaLXODR3a+rGyoy0Dg4mFHlYgVzfKM/r9zT6S
IRSm2+wylq1EWeo47TlM1ZwPcX5o/sicHRanvbHju3BkGF5NhLrMPynkqz+pvS4Q
UEhrj62GKaHQNKBIQKD4HbIEeqStwSMvl86t0iYIq3ta6GQAgh6n3Yo1DkFLpeD4
cPOO1zJetSrxkSuchT39qH5QiBhVi2Zy0f+92GkbOCSdaF6NcEdJ25k4Lr926wJk
z3fBAClDnjAoWxeABCRsp06L6451Pa/WpjEaTWWcNkFkUaF30n7CZ3I4TPEyj04j
O3h3c6KRr5RP4n/dOzkuMOyL3rIQiJO/tZRKpWAnvAklb9mJvkKcNe1rmTzepHUr
uQHSGzStxO/50uHcyvU68f3pwDy0Nr2dZ1WRw0g7Cd069PDX79ceFidJoveUjns7
jpGAon/W6tZSYEpM49gZmI8Eq5ZAVqTTmmNSiSufihDnyEyzkrTOy8UrY0qhssBx
J8eqGqj9ySJFLHJ+aOsBCj4ClM192SN4ea2et/CWgEmsGVTJ00Llio38RXId5KEQ
A6XpSAkdRQzm2SopP+J6Q3EJhr2Z9qSt/iTL07EOJICC3V7nalFqE+7zz8YeyPjx
nHlUs9qWnIKP6LVWR8y1JldU4C7yBBtzncNg6NxjCPs1Cg6GGNK3zC/UorLXCtmG
Me3g7ZGbB8D33I0V6lmPzJrv4sYLsSCwvgXBLy/9CE2ufq6BWlFxwijA4AfZm3pk
3UmUjW5qceY0/KPWfXRw5nWz+1nW6fuarD7NaBoxtGnVeVNRfeUUFBuUVi7dVLNE
zv9xQYd5xcj6bwtlZMwrgwMU1UaTD+n9uE47EZAEgE3ml0RV0BdIJdyfSrJ/fs9/
BBSScWqZSSdMUYORBLXQ6hT9oInG2MurDoW4XotU/qrURfp2D0uIS3SJ3TIayUjy
VEwD8lSmylKr71JANZk1AeC+mQSDW2eJ6Pnd7xBbBC5hmjnE3hlWx+9nmxtPzAIt
YSORwdrVEoxZ3LctLSoXneAdummytN9v0uduhA1NJ25H+SKKVjS0EzfGZdkunBCO
2R0fZRk/RM4xHBjWM8gO4K96+kdP8cWOhx7dEoUFU0iHrVtHyP+qJ6588Uahirtb
JTW6PRI5awNxp6LFbv0qf/2yTj7/13Se7bvX5OebvEa8nbb7wC2qEVmzbcYzV6Qx
tuM/IjwFbFyk5U+TOmg3bWFkmzBDF8QIbYFlpDijVv1HRfIVfk4iV3KIoA5J9bjq
KN5GeuejFnEtumSnMX0AhxF7u9sMt48+u1CnE4+z/ZZ9zu93lsPlQtbqTPsvmoH0
XmPQqYkQ6BxVw2MtXw4kbDujw0vmSriHDr6lPMjHTNyDkv6TPx36UvJyLsFOjq8v
XxMUmY51XKmduFUjXWjqqa48jXqLnuCAlG0x0eMxQdw4Cm4/UcU1auD6BGQt4/Dy
tuduZikjj5KswajVq5X9BNFqRB4pmVBCXBBFGWMzvb7s9dLVcMcRo2WUTphxhv2H
tkGpQogvM8QmM5zUJRBCmCznjrmP+6zhlX6mmT5Q+f+ehLCXqe0r0UMJ+slW9wz+
fs7KcD9/nshoJgYH5IYaiDwOsrYrTldyb/iWTJftZIPXvVhmAxhIjTBmp0oi0F/G
I/18YHvARSzPX6OWBCTLwj7IaJdyozUNmoQ//gcClFLA8GReAHwDsxPWbRbBuz6P
Jxf3ClgSO5wdOBUzegXv339O3xHIVN3TUvdmayAUqgxpUuTdAlJipq5seL7Qw9v3
+SgJIGWj2vsPoYayZqXAxrqF1ZWuG5AuZF+YFtXUe6Dn315SXPvadsLH4HYIX5D9
LHHAy1ZdzfYGvAmhz5dsvuo0RfQKQ7Wh10oQVFOMmcmUKHoC0zmSKmG49Vv9ezwN
qTMEBskvoNpFaGzsdEi1myqRNIGAlCxhSyEKZSfEj3vFchwEy0E6lcgCgwICb5v+
f9wquebtLxnvK/0BHJV+IuEnmOiqYBLEplcLqVR0lHQpnjhF6Jbe+cW5eTREgQQ0
RWXaYmNtd1ttzaoJsvPAsppDILMH7So8bJG/UHK+6KaHIrts60T7WypFDjagq4uB
2Txn8KUn/h/Ewu5QFgEM2LI8rYr3Fkm3czOMv84WkkIuV8TQ4+k124PK8J7C0hKy
ah09Rg+LDiVJfGFNiShGGOVvc+EsCST24by3SnCuL3+rniVpFe45dYgjiDzmoWhE
F4OlneRqzIKJg5ABvQgWA0SUQljAfdS+ZaG6dMXQ5Lu/B5oRI0b0biT82nS7pXjA
CVHNce1ZgGaStsaPq4rocuVu2jwr0qf2eR5aEV3zUDOnnNjw2cnGqKtOgIk/dJjj
lL0wkeyxaQeUaRGGITzWiJONH/hFg7lyyJhxr5+Ir13dRrbLt4qD7jHp3zDwCbuo
WM4dqO/VTBFnuGp9pX3DQxih+4qKvaQOhC6kcuLauMBPYYHQS6Jej45dJXBXEw6k
P0TlymH56+56GZfgJ5TQsS11ocWVT79SoFrx+/4QkASxz+F5WG/wEB2lnVUGioPu
REIvIaJaX8clAlhNUsuFawEL8l5I1B71IPsXNe53loLPndigYf1liCPTxFwKZstL
otuX3pARDZUqC9unT+EEkzlQ+XIRHW2WOecQ4Wq3GwxfWrbQ2jIFXaYWvQ7tiNQC
If1P8UK+XyRjJ0OjJL50cTOPHkjhKwygkuN2lZhRWYfCudmhP2+8kCNDdjDT26Ze
Ebx6cRyHblYCU6kEqznu72BVQoOCZUp14yDYMzSB8S9YB/hb2gEhGr8cThA09LnZ
044/A0h7CfIubltNXX5QC8TM+UZkk05NjGOlMDPlY2qkyfltbrHzOOJ0OExx798N
Xsc42UxNs14Ckra4+Apk+lbsPwVmJFmlzA94AYzYa245AeIXcOqDVf7ghdbonH2y
66T3el8vHCftAL/j2eVPrGYi/YDDKkUbB7uvInkCrcigfozHCCFkpM9yCIu4bTDK
8a/xfokyCP5Cw8EUMFPT7tUxA8bJbqQ1vrDsr5x40K24hbHQb4ZVvpQC7gfnTNT0
hf/s1sqs2gZQfvG55PGAFacvr5Lz+U0xNQkJ99+OmvI3JuhT1t0BUHzoJa3GD87O
aFsocEu0AMcSCp2SMSl/W3T4c8UTsCltkBEq/Vkxf6+PV0cfauhSeie/FktFxaK9
DepTSxGW63Y2NmfpZg2thdnbmDw/mWbhSAGxBdrzT5d9uVtAeRO2lWt3UfHkBqER
DbxQXyJZMpWkN6UoIevuv6ahVE0Q7YfjDt/adcOn+rvrWdDsKUtDUd5EUNhs13lJ
9zMI8JeUxYBvBjfIhurHNlMGAjBbc6+8p0Kdv1bcn0317hA7YicneCnSR6arqQZw
oQxNdwwdOwo4nQMj7U9018S/7QTf7CUJ+8O1XWRRmWfB2TE7ijEn5tvl8+Q6eduM
Z6BHbILOBqn9o3olmIYUCBQINOQA3atNc3LYCAG8WRxIjICbau8WCNx4nwP6x4fK
DII+fcfInuFRSfgY8cD0GkImtL8KyRayfz4x0zuT2FnFsHSSIKMpwOzA5zX3ntAx
mM1sol4gTix8+92l8MS/Qqr1IXz65xVyh9MNGbCfZ2dzYdTYRYltphO6CIydDQ1C
YRb5JZEHa6FMRS9/MA+/kpellQ0kAweukknsKE4pzWvRLunDQEUaJaLzJ817uo1u
HIH1ZeTSKu6974+UrcjZss7Z1R3M0HqQBQ9omGXmgIoRjZIhO0OU1z9P68v4eBt6
4V/PuQSrRW0vmIyfMNiyNHr73d5j+Q5aUT8pmaeXClXBNnmQ9tWy3w4pWLrrUCsB
holI/vnXpqkwHOrb/JpW/Q6AlfLSO8A/IZGj6j9ETbnE+S8KKen9tAqp01ES5lZY
Gvpr6V4Sm5KTijQuycwYQg721u0qlqABag2HVF4ysBP1OLHnrexSTv0g2iqZaAgZ
5E3F0ODSnn3jGJUEoMugwdJUMamcjzhn36jjqsBXKrkJHMHlFESp0RrX+9fIxLfp
zezWKkTBXnStLBsAbu91WmTOPxjPpz+Z/ZgiamMqwY3grdHsdmmLvWUWiI/HuO5M
G/HGE/ptZjaPebq1Kf6eTWtgwBtKEsnicJIDJxaQxjkVQy6Lcv0zOSnKigq/ENnv
7ehBp+ptzz9DRuHJPhwniU7Tfmu1Unkf2/UefqXyoTqRm9n9R14xPGcnqU60uJlJ
CLk8FvO20jaYtUcYns0AUYBfXryKGCcuJWitIbWlySfUSX5MkgY+5HZFEt0uXLBV
/fwMdhJtdN4QUre6e5Kw5GJLglYmr1vsL2GmQ+sNlr+qCjOJzI6yavCczkOwKAz9
50d8tm89htxrnazCsCRBGkH/SE2meQgBMIPlwLDM8w3WbQNujAdgxrMj8q5ic57c
GsGOKKlTArRmeHNHiMQfLj/9Vxc0X+S6B5FlVg/b5ZoyWnqe7Cy3GWIhsWz3yZ7P
Cq1WdCkDHF3S5a3Loce8jbbsAJNh58Klx9NCDA6hWnrE+qj2yGWFis6PNffFqjd7
KNDfV2+en73GrOPzgbjfujLm4fOl13wWI8XizjdacGNgF7mBhrLwv+JpK5zcvVNR
C1k5BqwFftzjpHQTpAHOGK1wT4AKIXgmx0E9gKWdaXqP0rb96c76is/DbfWmdHzF
Ju3zBXhcxaSFVYEf3rBdiQgbX0PyPbKiLTb70tGJJzC7zH+lArPH7FD0t0+DzQNb
Ibo7cAichCxgYzaVXVkOBeVPlPm/VoeY1lYlng5SJI+2ReclWR0ZfhHo+0UQtj/A
o13WSZJOC4GxFtQzB+DfQrullRDxwTDE9a1g9dPDpmyLbUMjNCApOcbnGHI2Aoza
GsKoLIRykR2EuQFjaojvETTGzuOKCSrgeZ1pAwr9UsOni2KIOFE23GYva39RdyZv
tNiLlwj8fuJA4oW5lz8Uf/RPNR6vmFujNB84GVsa+vp/ZqjVyDQdUQHfUAiaBSNt
qpUTIlja1anPwYvBDICCIthCRoGxtYABawspww9e78VLuBxJzPtpcyNh9m1dd3UG
UVXCsl+EwJeAUeFUc9362ZkTs28gV7MXuWyOTnoxRHolt46Dmct/5wFXC+lwBluf
1zia+6moBpw8kaH97z753rhYyYaCdqqpnzlxc93KpRGlMxIyNVQPL/ac71QUVXZg
9OPwpnyC+f1eie50I548+QbzakFW4MKyuHR1H0rmneR8cM6xmHBBUJXlvHHRPno0
bQEh6tLAQtrJUejmWf3F4QbCHwmZFFtUBiljgHfS4HDBt7Gp6W4Iz2NwiSweeHHe
PDQjdnouRjLDWTh2hWslSjejkFF5v4eshsrNfZh/voxlz56Ku44MePYhKpmzO0b3
VP90U+KJZ7l5D4ozlBJgljwCagbVm/YhXI3Ba29VJtVanlaUPGF9bbAaD1KZFXzw
nny8Pgn4RdHfGn9Ogyf2CIxprGDnDSBcJYBI3ocGQKk2A5iCmtuMuGrHuPuYhfdX
f1XGxUiGKlE2+wx2dce03G6cEt7FRYXopWG21DUIy2q6W7FVVHrl5DTIod3YOpqS
5WZSnq3UufvinXIumbc2vNO2qO9UYeiopqVH6nDd+NMTY7dEQpgWsdLkbksEFY92
VK/V/pc7N96LSu9CqjJOV4FjXdZd3rgZHJ7Prk7Zs4ZchFthcf9x0a+nVrlFGLCP
8vWgqViLUftCM1BYe0t2vjG6fLJnvUZBIw8YdhkSHxTnrblMtcWea1oi2o7QffG3
MWP2BlpOBEvJt8SyA8gDkJNNpSgs1Ff2uxCKp7BtdMfsaPQbeFy33PE6PGerngqv
V0oUWKvVz3zb127/MV10gWrw1W8Ql55eGdQG1E9Hal0FXZCRuU42kT4rhcUnLMkr
TwijMRZMWpbnHNYYGptXFiRP0P3an/bbdK/OnuKo+eHbB2YyogKe+adHw5XbVWpv
stqMomXti2r3YZvdZmo7zKWLEs8+lMOvaO7j9cB/oOs4yrPyIB/PDLJLo+Lvt+3k
kP8/yeTTSwN+BtFivXLRCRlkrZugX4qTh2oNzLZR9oFuTVngRTjWEUES7Wkt2Xmq
iuDoh1TsQoVB1Z6jrwC+03stHuufwIMxK60/bnz/Tf4MCUPAOxAj1r64181lc5sN
j20a4dtxLgP5bEV6g/9Ngm9kPgDyf5tqjql/tb6A6qy4LhIsAoLvj4aN/UgEgQQt
qnpIJHCdNE1Zj0p/AWgzHK6zo6/23Aj0dP8fVyHZUwbqFx48PJ8iwHaiBXCFpV9A
tHZcUW+D5xQSRR8b4OFn0t1TdMbxHEOWnxhENDRwBEaaJlzVPs7kLFg4HOk+r1N2
bmOJeADoex9BCbDLnUS8IoG0JbU+AB6r+JgRApLo715yqCmKJG/4+dsN5ALQhU2g
IW0ZLLimYGd/pHwu7xzw7QMcax4iFBoKAsjAYHkPcg8bkWpb+Z+SPxpfe+xjtoMW
VOwC/PitX4CZugAYseezBlP/CbXX9lPKlj+IrztLZyghJJDHFpsA5E9Yjq590EDs
BsfSMz/UAdfMyJ0nJ4PvvSUGbNKX13i/IrCY3XZg+BndHKefyyp1xJeVn9CT3JOf
Rz/O+K5BOYDiI3swSQEljsMAHF/jZ+WjEJwvB6XtO5dVEAU16F94ZDwRd9C+6dMB
m8EOX0ZlVakNE1qhvLx43s1opZSXb54YOJhvkMLiTbieCt1eDqSOP7gNgKYDzFzp
UBSNXUZPQtOKIrG2LPZndiZdENfdgsfDsClV8vqACuJAv1uTE8AMBgLFzFwx3UMk
K7RmpFFgqWN9JnB6i1btSRkBTBJlo5lyStbV5f8TU76KHb+DEp5hgFlYKaRiHMkt
zw2xYyoLbeLog+B0/lvMYZJF6D7IP74eb0WeS+rWGB8TFicXWL3IMzH1tsQpU0eq
VTvthP4vdcefxqbmb27V2HdneaMKRtkFh0/9uq0ZrmA7qQQ+lWJA7EHpojKwLn36
vdQa7bIxho23NLG3cdGj+lGmAMe2gCWSX/xrhtkcz3q4f2KWa4WSv31/j6TckdCC
mcWTQU1YuP6YAV06jjHCcenHQgd0qY4KZXbFPjsDh1D1uj4/+z+kOPl3E54eMt7l
CcDSRHI0eZEl1/Xf+UTee8VSOVnBFEoJKPgzcStWARLtck/yV1i/hjrsECNVAsPE
ySsdaoZasGfisdxWt4U5/8vvaULbYvsYlEiVijXQb41zFncOwKCmf9QljFoTepNy
qcoYCtRdoFVHzQ1NIzgusm5BhWaol+kfczL6caC1gGdbnwK4325NolfxpvwOtSiv
n5/WBQViB2OoMfq8Jbh9Rb3aIqc7J9xUbR69BuWBH82IME/f4AYSKnUfGUSdEj77
R9eBSvMhFTvW9d02pRp0z5BN/16ldpIE5jBV+Gm3jY5SLoWL/GWWK+Qo1aWgF+ml
dTQHkli8bbHo2GPKZw2yjehd1k7rTQkrNwcjWXscq6j8InmEtA6quq+ZMtgq8TXT
Kw4i9OiGbV2JuuBx9w6nnv/Qkub1w7xC3tDDi+lOZm3JMHEcF6aIg2oh04y3QaGO
ZddtCk/yJfv9Oapj+vpLwVkNeodnhsl1EatgShsuvw0mVwh6sHbKjgNlyRHSrhPk
/zbKIjrVWj7fLWztQSaaKlndpz/jMf9TT1SQ+Gj2bg6lPmc12jM3M1l9SI1CjJ01
bsv4TYeNwrqU8Vm1z+dtak6FNMe7/J4hGd4MH2bjNeeM+m0lQcE3FEd213oMCDQv
SvfUgGRGgOgiV+whbUJDs+TlYS0eDxtndEPSMOmHgCDxEuj1JlGhzuw3whT9uSi/
3Dcb5nCIxb7aVIrvxh2iwhlytXwPVrh3N5nvOMJUPbGdImxrv7vP6lrKLTqbywhH
8+++Owb5BR5GtvTDUDmbTG3O5+uXM0baRpbTsuqzplubioKsHjszdpA0kieuKrtx
UeoVMpCS4iklPFgeBuvAp01ixQDGDg+OpHi24AsEe+UhpFgv6ZL+PfpHw/ienFYO
V7BiCuDUgTJhdYnsHSclalYbKRtBevZUonirEHPFU/uYeRokQTe1XMUisKCS19Dh
2NZBfsMVk3s933/5yDDUi3j8QYkqPOEuXQHdfr98THjem+xL1q+Bupk0k3yDhrLk
35tb4fLJMpNwlFvgM+QOOfmKGiQPkg2r3sAPBFCN3YTdGXvke4iRGiSaMZEKb2Za
QFB84/A1sAFXI7mav2/KuxHdwh+arGBJFpPb4sB8PhIYh/cL/zUOlyrsJaVypZIe
jglxwZImwn/uPZqDVHfqKhIYPs4k+c+5gZFkneJ2ugLoaCn3BYeixYdiX7APG30I
6BOYiCFKaXPkL6Y8pHP4s1/+YrZh13minkmKm1W0rJs4rmWeDCOFcepswlO9CzMJ
OE7pfX6KxUdc6F8C+BLTPZLnKe0kNi8ijoJILb/I03n+4Fe6AacAEsKAfi/26K9Y
T8vaPrGT9+0W8vAr9TYXby/I7vkeVwC++zN1lnn3PIff1bu4aYdR+L/DS9+WX47W
/2cwPKZs0Fgui6Qc7KlV36J4cvEAuax4aMy09nfGC0Cb0X/jqM/8qOK1Uqvn0Wva
FmGopqH24MHhgyCxdmkQ2kiWqR0zwX3ygMAUxAaz3iK9wwnGLmehoLh6ZNhrMJqs
drmws0w0jxu24fu92mwfEBbJqreTVvH9rJnUVbemTQ+v6b/qBDg1KXd++T+maKuc
E4g3lizHpKcr8SM+s+xcUyAE2exriJ/XzQsfZe+lCMV46clL013EeZSxsC1lkw3Y
/dvGgqEhtdoqfLeOsFhBJxwnBSyNfAQd7ogy3H/dUA0bBrVpIInpdXH17VIdbaNn
LrgYWgdiKH3d19T40j+ahirmnfJFSsRE56lcyEBvWLgPNw4rc7nIJ/rNnRo7xj3+
bz8ZqClNsRCtAhl98duO11f2zWAmdN7PUWAd7P293zghdEM/XNlY3i8joJi5yr2E
2wMbVxLva/pxkyyFHRCTMyujX+T8u/KpkShhjoYRryiFZJFOT1wUNmJXrph/hp6H
/mN8YfMXNtMUsfilmEADySyArQpQz9yiUjmOsuulLWIJAjCsVT22BCSfV5ztfwGk
txGOdh9XwQZyRUbtrfsMZGHuFh3CiY1HRmq04PKXKdXaVjW7QI0mbkHVVAPLZ7cS
wNv0I5xlSmE7HPZF+aE6JRDzWe0FeEFl42HZAtBd9Jn1ZnDnU+RYorpTZIag3hbp
A8jaNg8fHuv/DK1jctkgatFnE/mWeXHGJ8Kh61FLs5pAkaRqdjOVqxPXZNuFZ7Ec
dR2czLvpbF1u8oql1Teu4WY5+YwKXHo+viJ+LsLVtxc5jtTngm+vxmI/vwCdY1od
a9MC9DD9Fdw5frvrS1aBcIH4eLNg+FUnNIt/Vhb/pfo2S/ZFL/lDM9itzQhNB6l5
K1b33pJ1cxQC+9v2tug+Kf9QeSPdKYNlRvzJhpT18+naTovFPB5oXlOBVbmJVmNt
0vjDUfIljjoIVh4zFde1nqYzEJhttwW0mNBh6/jMV/L93LND6GSkqjvuIh66NSQv
+aBqtw28HcSrte+k/19BpKxFrayR2SX2DpV8nfX1jg3Xk80ErK7OQ4RxW/YUBsLL
smRoqDoaecxEJMgIjJwv49f0rUPXGQK8hlLWB5FZJbqKbZm0XGpMogC53Sk/RQXK
gy97PWysPe5au6KHvhqimEwQeSGpR6GkSXIEWyXKzJFvv8exuEC9x/VuLveHcsJF
eW+wwqwXPAiW0xTpNapCVXPDiQ6T9FSCwuF3XwCCIX8cHj8O77tvUSWLEpzzNOHN
coz1gw+ReBxIE8yfmBkQaQ408gqZHsT5XJq5t669W9lvTGJIsufB1fLU0zFsk9ii
iKQQ0Y4+DazopY97d92lcTFEba/o4Yo9248LSGb48/YjHZ0Am6Z4O/8+e0IjsVj1
6UBYY12hSXpBGBkXznwgqUuSctpgXI2Y3fC6zz3+FXu0I9+8sNr7ucWwauJexxQ/
+dRUYsMh6AsLwcJPzkWl7ql9sTNBWjVZpDzHsyPDmkQnzgKo/Wq4/ADoOgFmTu9O
R4nLE8qUrZ3j2ffKcrLFJwk8bHEEck7oaIAIplsCjOz6c96HEqw5uRCFkmJVre2A
N2UGNLTLxzKEHf2WqZkMKiMe0/CnwH2aU5Tp7eI65ahTx2HplB1OSi3iV3OEMqk6
eoVmGCaTJ1439WZstKmQxQGI5iWttC0Z9u4eM2o+oaTB2LtZB+wSuZQkl3PaNpy9
t/FcdJBPz8Sj4MxPf+TXr9zJ1rpOn+uo9hyoJl398GlkvdZ900quUiwjRMLfPdsv
Qm1LJmZLNIM3MocBKCm+gR5l+zTjMMQCezjli8QITVuupE4Ugf2WagmNFh1bR+Z0
J5dDd4MBk003lPPf2GPzb/R3kmdyOVZgtLhDdY0PAR1e3iVKTBPsoS/X4uhvNfg2
bpOIN6s457SHklLf9UuM8+Wn5O3H0rQxABxa0JV9ddIEHL2lG74aGWETrwzQWKxq
Hm49WFSHyvuBQ0fXPKbnl4+6FSm929sAXjznAvE3dkMp5uVirHYX6P81NIngE7C0
b2a5DOW3o2ScQrgnp9+2FPShTcTLyCMWECr6ShFwQRhidY5cpb+NUOfVg+RLnqbg
U7qJk/E0SNSwFvhbvxaSQGq31R3sVI8o8XWPvSuwyAnXUpThed/FGnnEQ81tXdzi
n+5kqYQ2U8F9pjsLYfbbAdyynq7J15nFvDYqxmpFn3vq6jeGpxGRjKQvt5UaPt/o
GASrm+Q3CIH3FpPfbotE+dKNatOEVBZk3OzJrKi6moPn3x3r2DHabIK1zi6eMZIi
CX6djPxMlfytGLS4SFQ6Klbh8LdsqbDCWkE7+unbvGVGs0EEhD+sQFQL+28o6DdG
mislTlWPM49umcwGQqCtRCvlodiB5VSzUERcUyDv+2TeWnenD8JHBuRzOV3K1/q/
g6JmNvTIDCwdLaTxcY3z4D+CBGwM1sVkHlzYNiacuBONvUP2BSzKpPUUxrCivFmN
0Xi6dcdhuYUfM4uSf0fqmI1CGOyOwtWWjOEtCqTeVXuBqLibK7UnIga56b/XOlDn
ud4/e5Zbz4nBGhVkGpqZ05g7q8VfDrxxAnoVRiOdMHF3FNZCKoXkrt/ZM5DHKs99
W72zeHadiM2RHtzVaawTFYZd124xriUVqG3vnINmcZjxPzbCZaPP8Ht6eOhpohs0
9ErAokzHlQBkbAju/CBORo8Vr05Rh0lsLCLv/qwCaopQmrAhUPZ7RM74uXaD+Q/f
eVIEQw1hh+dA1AZ2I+JcVYQaBgJl+BlIDSMx5ZwI2sxQPt38hakTvlwTO7stgNfq
8yoEZMBnJSy3Fm8r4vsdblZjef/kkQ9u+RBUOrsk0rcCLJoChcfVNAo/udi/qJCy
LNob9dMZDbkTOhWDequjBea43meCuYGdGb/b2JJIzT1XnK23sdySkvhaUxscH0wD
FhoS/9YhaBCSiad2qRTbRb+fPeA8EF3KU+7A3NHe5tkbQxpxSfzPZSsCmw38gx3a
7LY46XjVUyr3x0772ixavm/ab2llgMioaBUE2rqqypxDBMumJ3/WPavhOFgziHfU
fHFVNfY7K8EbxWOGgh2+SCOH7Fp1jPNCSBIbkPQbMZFPE+ss7tmGft6jvQIdcxr7
hAXqVxxnyk1P5Ko0xNURu/m9Wp1XxErEqNR9d7nGBRZqUSATXDqvZkCZVwhSZh6i
3h9n3JRz+rVpL2rjZ31wtkn/CQfbp+rFh8c6EXr5+0DpSZt6HUICzKuKkqX7az0y
KJkmOv+ofS/RiIn89MwAUu3frEEPm+kQ+U8vMx0R6yI3Eex+EE9Hsxo4AfV44Yd/
S80yDtkobnCmq6TKbdqOvz4AdvEb+ZLU/YhSVGkvacpsomy06wAYHl9wwRb3W4Vk
BYPN8kKZNSEyod2Cx7gRjYKnKCjfiFspPV2XbKD9cyIx7DOennDl+QSzJ/sAMYcC
eLlycCMrVNQf++8O5r1SAQAJEf9H6l5hkA+bJAcOpPJb1pgaF1rrUwpDDwNtZ6Hm
qSFGOZeCNq0/SopYLBLvWG5qcaISJ+V+rlDUJJqNiVcSso9oOeE7fKmUiZ1GWmJZ
NxAy9PYkDoYURzW/DLf4MY9kHp1rbng7QIu5aX813q2uOmroNPj4/7sz6OK8dW1S
ilv0EiHz5WB+vVLbJA6swtu9yS0J8H1ld9u6cQlM0IZDqBJulINdGxBOKMlTJyl8
E/zowWKwttPBi7OgU0Bj7jXyZAiQtJUxDtZa7pM8F18Dc1PXgDvFqhSFWw/HczYL
FK0ze3wRQ0v9y1dwKmUDlJFTVDtancPnGlixahc1BgoOmYP1/hQRMYeo4pho5yna
kt1RbsS8U0OOSxnHws7XBnc++lu/nkaRlzCZhRuP1Oe5efnNICdP2PmTzOkQAF0S
D0ewot7z6lzwvQ2paJDkvd2Ssf+uHVxYSGiOToTH1p9qSOkvcavcCeI+DatrI8gP
llSWr7hZBBq8HzfMOpjH+O0Vsf73c0B6+xQx4oJDM5kadZW3tIkmD8OCaTcNY8SZ
nGQyyQtsGgJcicaSw5R4OeF6qDdsgKkNcWRTIhxw4/7CVPkakuYCZL3veNMbdG55
YpkaIKQA9ByT0StCGUE0Rq9Nn0Ty9buQ8LFeI3oGyGqGgnelus/P0t3CR1WL8tTs
Q9sRFRJqBMdo0oDpXw8mgt/czpZrqikcGTqQy/5m+ish2RCX4GkzSiCCFySLe87N
mGC5H9kQFBmxGi1gIJFlCZ20CzerSJ7XcvjZAVlTaMz9L1pdcXHO/xMF5cEB9YD7
OxfRxn1HplBXUGTFWjiOOqkeQFW1qWTwa/DcJNgtAGnH5GAWbXHFrGl7ErdNSxEj
SzwfLAVYHXil6IaeVvdpxx0omF1vSahCJCAb46o1DdxWIMToBwAUCF+cGu1xlsiy
tlXpVdO80oWp9BJSApF0/1jmDaZBU036YE7ISzH9C6W88cacaXZi12tCVZW30iNu
tFWPilurPRD+T92BYVspCRcUWXndfQ2msq78y4F1lHI/d+gEKqh9C7nHBxYCAxMR
dM8P1rdjnSBxGFP2xwHVpcI2qIC+lyis+wmvknpRq31S7Ze8M/VLK338EIZu/qD5
9ftU0AYwVhVpg/qeXXyLKP8f3PAU+cEwL69r8rpRB5dASjsU/NoKK3zgI/QDUsyn
K3dlD3GnGWePqgIH+YaCTO3WTTCh/gUYGsxLkgedYdJJBjp89w93cfJyoNdfAGnI
fK/GX0whJ+otKEef17SNO7EhGOv+osd9SN9S/sUjIKw7K5ltvk5MiKiRFTD1NmgB
xMwKqW66eXBea4+ZLXi+lKxWwgeM7+3TctYU7q4POeHcB9x5yumDeVRb4QApDY6n
9Ecp+68NrVl824HnM0D1f/I82dUo+a1jfXPr2ZQ5GjpMkyWUxfPyW/GtvyePIEHG
nP+Np25HeHnx6AKKz/8JH09fzrafa3KTKLpmb8d3o3FeOOmjSM9fFYGSS2RVsCAI
lgJdmeKBYnFJR0swgO+6fjktqK1Y9OVN2z5Bh7P2OgyMwsMZ4rBSQmR7hvWhKZqN
gK+hpwX06nNDmxcFKdJNjBi/wU1X6LOqsfColY2Pkfitr26G9YY6xNzSq6CtWyxN
tKj25EiqVmLK3z8v4j0XeCAqJQETpdBFYdQ56uJLJWGkGfCInlFE0a4aT+lgOXPE
Q1VF9NQkNkgdVJNpPnwMDska9JtKewKHBlsa4yJYn2bMgVp4jw7KFP40wukvFww7
It95UH1JGWuQDsq+GgZlwJXV4mzrXDRSrolC892PE5o8seEQGygLL0ihaSjTGSqx
Mlc/Aok45/yGAlbxnoBgVhpVcvJOlYy2yysxhnUxqIFOufI2Na3FY+3tGsT8/drZ
omJ2tlQQiutAPJM+y6DDs/rtc+M3CesVsN2thxj9l624H3lNNooTBhhrT1dd9f/K
Hn/s2l6E94XaNPl7Ld/IxYHBTjs4z/V0PPHw6KPNFpjvXFmUlaYv7PzPcZaIY3pS
a/JKrvVBuW6hnABfgytf/MH0bwZlnpiL8ODnVwWY0fCi554+LGREenR8bMkiftFA
sUkrWbavod1I1Guxk4OCIOApxY5PD25BHwf4wXAsGTb9g82gMQGdPKMRQtXTS9+x
1TDirJoMcHmxJti9RtLFcnkDKuQK4/auFtgDg50pLucXp4slEQKvU6CU6cu7nq3/
LDtu41zvac3L0aErbxIxNdwHVMjU4XgHJpS0vVRCY5NwWzrzS6IFSnAhPRuZNvuP
uytVl58oCpiC3kkY1Xn2JVvTrHNpBo35qsoZ+eu81yNrLjZitSsuliq7hJOULg/w
MiWrB3JTcRjsT7HuYSHYPkTt2lBPLz5l2YgxzqQdd7kg7bSl6QRwgqTv91gZDz39
jivsI/eiUhqW6WMc9g5GL+VA+CB+5i2zEk6nFnxkEGXg9HpBZgnpHhJylhlfu7w3
aaHx8/d3vmrfBG0VxaXnmi8NkiRNsLnq1QnjInEOZZ9Hh3jvTOHJ7xURBifKz8Sm
m8XBllk8i9L1h/Lmudyh2H0ForRHFJV0djkPVloMrJyhClMaBcdXDbbDkjaoZX0R
ojGwqt2T2LYfcCRIVG2934mE0G2w1N0W5BzarfJHWDCPrGosYSYQVDLlkxWlRNoE
px7hER9jPFXxKVh+YqgavgDfhTlgZ/wWi7aiT470KCGj/SUpAY2upjFnB0lQGwr5
ax3L42RSB/DBA7lTmCscQURkPqAZIezkwvFD7Yl3lHutEFSP88ZWjgTLHsr9qfam
f3P0X4puOZgl9fd2oIQHWK3E/fNpor+c53UtI2f6r4yV9j4G81S2/urtPOUkg/v8
nw1A/AZ6OKLD+VgbiYe8qcTBtHfjTMSibdBPAf5mWOIH1EdKG3KrwgKprJOlqtU4
QJJH0Ei4HWNvcXIRZa28jkdsD2dNhPU+dKO4oJigZbMJ/QQw7lgIBGHPAlMy0U+D
ys0fwEex2mRmZAeHAUvTC08EeBx0OmgCnwXqN3GIcUTECjf0Mx9biT/rwHAGsvn+
HIZiND1Numn/0j7s7+T7eQ11EeRvYCFVejrHFMevDcmlozzkAaDdm+RdmkXL/xAV
w26NwA2iNnTRgZ+cVkACZLStgd2Gabu9x6VLkyoyWLxJ/LGktXpV0zlEk4Tx8PKd
Jw16tdWcK9Tzox6huGliOXUw5c8Ts7R5qK4kpaQ0JRe61LwSQVWZDfUEqB2Ty16n
uYg0S9T/VQBFjlxtGh/CWnnhYC4/gyMpE8Rjyt8rIVVH6D3DPzTbBLWKemRbcu2s
jrTlJifwRAhoslFd649/UVAgJrn9IFxbOBIGzhFbbaeX7eP0MBSd0ZZvFhQnfBaO
AM5wgLtWTl28QJZWUSURjlu3Dq4yYuer0bUAgWoixuZ5zUkHlNOteC/XeTu6CT8r
KFF5ySHFuJJ+rlmIv95SHgS+8GkfjImF2kKQj3RlmK3jAdNDrUctY16Rrfa30fIP
Sj8eBQLbUasKCUvpOp68FLYyD/eTU9ZV9VNoiIZiYkcSuj5zEg4Rx8e03SDaLxqW
MDOmjJmb5CzZ40FPpJfQpGQWfUOaU+mdc4Xgbg5/onRA7eIvsvz5OjV1qeO2h073
dTtCrisSbS6Ipl75StAn0M2v2Ahxx/JN/9sJ6SFetZ9cRtz4gVM7RNyaeds+GMMR
fz6NdPKzDgVaKLJPTo5AOVe3vdTvAuh5WV5GEPGmV7Rfq2BhtoD1vDfcQ9weGGJH
gNVFNzm3gXuj5A8A/C5kIKQK8I7R4Ex47km7HbPlo3xtZYyBMaSBcuPIV3tGtc7t
/YzwCNrePIv/FTZDXJZFn1W86RqUhHrNOCeBc1YRhrZ6QjuRD5v+iaXq2048FLP9
SPYX1Zt8zlm+3cXHzGmRQeIyrIzkUhyBaiu/zT1edHCrKgloGveYPS0F1m7EQX+v
KNBevZzfArMzQCLxCkKZyH5UNvq6twC/TOWEFH9xy40eZEsFoaIxes0uaSpr7xnZ
X7jLK1NxQ7tQyXhqZy4RAk7CI9yITKDOIGLzxhx6kTv+HcT2ixXcoY7gIBdaBSKM
GdMi8On+xXu5XflPj6g99EW5d1adrzpakZ7fOCnvAyA5fb4TJu3bim9MfIpbJecq
AhLN1vo/uqhkHS7nVLMP1IXJe2u4HmV3UxnTNr8u42Xdyw4InKCz54WQMQx7mRYj
91YvPhSbYcRNNUrn1fmBYzNlpn7nl7F6FZI61+GdoNEpIyZuXclZ+/EI4ZoxKYRV
Dv6wru2d4udGPAGwFMKuebC6BuKDVH3dBqBn9MfYFsd+30Ct+/WuRYh0L7P94VQd
UVGvsBfU51EYpHVmP0QrjDfW4vQfIp8khH+syOfydx+Jf6BRUjd/uw3XZR+L3BXY
c8dttAttOtNY1MmudRmnHvMRL0yO0fS1SxfWtrIDN22H8R1hDTT4/jb0wCJSimhw
KijQwDVbf0QlvMlfFwgX03EnNjvajMDRLD/NIq02hdUBbY6QqpSm12klnz7urbdw
1ERGllk64UmfYC0cIvglTfZRtVsUOJYVg5D6iKlA+7ajCWD5EVKnUtbnJVnrtqct
DQ3J3z+UXuiCmVXvMHz4Pi7IjAH4tJ0fVlWbZXZPrrIyQcvUf68CsMR+nlr2FgHC
03LwgIRlOxPbFYOK8/rV+4mgKeyHciof0bOPNJ85+ao0ln6UZ3hzeD+nIfV4u7Zn
87oMVOw0kvtgyndykSLwFYFHyDdNqt3uDjn4I/DHaYQ1rG8H4LvgTYUrTfkx80mM
IYGLsNo1pUU5ywNyV12EmOaJQNpjA/bTGLn5akvX829ZbmsSgPSYCUnVeMw4RNf0
wnK/V6KqGIsGEXQcpjtqykAe9Tpmsx+fWA1bHXlaB9Owuw3ElO9S5XizakKLbeFD
/SOxiuWlLGMBeqkTwny7aAL/Q0JmRxKrLjYzvsEpSFALbQEfRMy+5irjHoIDQHne
JAwreiXcIskaY0c0MSHzEj6x3eaVRxTi8IFB79MqbemRHLdrpVAAOw8bsd10d+6z
t87oOSzZb4JNK4FQOk9ivjO/t1XF719gK0G9x0gz2d37bxDuLHY3wvJQKIRuk+4v
EZD7TAvayihChW702SzDE8mSekS9JU3C7d9Nk0K7/ZARM3XdkfU/e62+cH2Gr+Dy
/0J3PSmjMO4XSALYEG1eSew2Lj585tjIhvclBeDyAwUYrdM5rahNFZsh2DSYxWsZ
vSfF/SzdMfk5336L6XJ5NkHuAHEgr61b0hsVP7qkaNgifN/rt4n5wBor7jwyQnDr
6RgFVru31Q06A0fZsiaVAjWLXzf+cf8Qs9hI0W1enK6BemxYSOY/42a7MCcZjVub
CqwyEW0TkhZCR8lIi/9O5WMCPtCjNVHxTiDM2AXGWdFn3btA4P08/iLqIC96n5LP
phFOVW5X0bIbuleCosiVY7D6EBFFvMgfFnpHXrfAlbgx4c6WZ1vlY2QbLsv9PUht
mWXZ0G+T4L+CRx7fht0QIDzCy8NzK/AxR3BgTqlm3M9zCoN05sHPI3H3splujVTB
qUTDxvD2DGYtZzXMye10BYl7hpqJQDh+MMoHJL8jngJSHZipjR9uWQwMwvuF/m4f
30Feye0PRmH2ihsmWN4uXDQrh0OpGqzdqId/hHduR3+xjfqT2r+RasvKoigRRZl+
+yJGCWmyQWfyo7+M1qlLVB9NOMyi1jYPzkxP6k2xA7Kv3FEdaBulQEim3GnJApyY
W8/qxDu/ccLSANVbb4Unw8fK9AQCc/K2nXkLb/DnA2Gke89Me+uXGpFovkoQZaya
7nqPU2vdXvaO0aCkuLH+8YTV95F1jVOL8g7NLxjQpSSimnz+/pz7CLyd21akX3fX
f/Dynm6GQyjbX1VOa9Y1QOkSGVRReROwz6L4P789oDNNJ/glvhBAQ4iichaJc/eC
NO7O6swE8nTR4K+GbXmd1Lr5LhddCkJvFin+6AfOKCkprkAzbwrHJZCtv13l8pQf
6kMW3FsCM5amofK2wB9vCKPftZxflEFIB5cqxp6+H0jm399gVBSnYC7EU8LgdR6/
XJq0hrHCQmLlgEn1FW6PBD9Tx1KWfWVmq+uZHXC45eopUhzTDUbWtLRTcSmIIkc1
EX64IoMAGDmeiyjPPmeGwoDJ2VhYuPAu6cL8NpCTQ+rVTVaY3EKkelfUcFKxN8JA
yj5mqP0yY3qNE9zaLEGoerakX9vH+H20OJ6/Cns09UNlgi5sFAnGeFrlyRKVPMJe
XxWgrVdZJk/+1TEkrZ2Mq1tN7qaLuj0Cu0/3nnDwhBEFlv/OCKE7od46IZxXCcm9
Vg1Ds226x0gXqSc8NjcHdQEDFrt3ebwPwz3QblqyboulxxqOsCyREVu1n4LmZt3M
OixNynkTtx83S1wy1P5EbJNDjC5RnGBYbZxdLjZ/ZXpiesE3zhYEvMmfKRpoZ4ub
yLDGfl2HfjeEbBfvzBNYbXSck2vXzdj87vfX8iJfoK0IfwytnW9+Re5IAJj5yoq9
vGFdFQ7zNL8r1mNAjaohRpB5JVjAywbT9jTTfzTGfIZXpZoxGWi8Q3QP09N+XZx+
MXgpjIK9uEaoTnoNuzkt3GlEPlG1NQVwHUvbwka3icMwbcLq6CCXXETF3p6b9Q/o
QLVGCLv9wFIL7gp6+/Wp/MVY2b9PB0NKsES70bLCn6iQpfqh02BLqn+qRItrl0qJ
lxsa7+fQdGTQlhv1HNuIhBkHJzoOXWKYJaeQIz5QsYP50bYHA8LZUUyhdKumI8pr
/0taQvMjj5w0NeYqCL0tRLekJg7ySiEayrwss9IdDXCdLNBcetaMUpB1Mo07ZjnX
xKTuAC9TdLeTCivL7HBFJsGFka9Tu76nSt31qFMgwM+JmCVmau++aF56NII1Pk3L
1eYjdyoW5yGugD9PDTWrlglaj1d2m4ki1SyrxiTk7dA=
//pragma protect end_data_block
//pragma protect digest_block
qK1OZ7iWJycGsUf4VzxaxSCHxT8=
//pragma protect end_digest_block
//pragma protect end_protected
