//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
EquBD74BMngxkxWqAC5LN61tNx/kfOxr3Mrt/jUx48X7tnZgI0YUY2glzhbZ5gJ4
2uDmy4KANTx8kic4V6iA663W7PvHlRuWtMOaj4bPWj207IxBdj5NmtJEhBoAMLGD
Z701OyeNZxxP5i4xXKJ+MQi9P+pk8sIyrEv3Nt1vwKfmE75yyQ27OtAa661NZve5
o7SkhlCCw8xVabfheD+uP1PiZj/2QfNRmCa3skAKFkhrOPkEXQ3HIKUhyp4g6Vuh
ZzLSJ9Mk97DK3iYOLOBezklLRygZBlXLbnC5lxszmbVWWovORMihbucUANHzyu4m
yXVtDFSg5Xz6FbVQMob4nw==
//pragma protect end_key_block
//pragma protect digest_block
hLZYC6o+rcTO3OQGTg0R3HluotU=
//pragma protect end_digest_block
//pragma protect data_block
F0/vMBlqWu44jbmRr4dujxdzaNephCa0vQGNTcPHByxBfGK4D8v9/YMnWBipgiiW
GnEaEXwtWQzhUUPN9loAiXaEeb69LqorTom2LuQ50FwUJHBM33a6o3Su0bG4iFhc
OHaMomSczOPdJpQ6PojgrFOWaIVmnaGWZtbKXKQI403yOWUk8mdH+QV4tzFZJPIO
svVmtFDhTbljoW39lI/zPA8lTq2I55tLmLSisCseY6j9HwKztVGprdkFZ4WTGLTX
BVjGGqknySWbk71BttZgFytI38uwzUhFxLGWlzmoGalN6Wkj3uA4H7uOcD804+BJ
eXgxphEta8UhUQ+iq+aZNVQ6BQlqtvDcLaEbDeiCEG1PJxJeKbzE5XwTyZiUlEza
//pragma protect end_data_block
//pragma protect digest_block
JfvS95cDbigk7fZ0KU/uH0sfyr4=
//pragma protect end_digest_block
//pragma protect end_protected
    `include "SS.sv"  
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
dQQ6pHjRhM9+xcbUwwj9LBXUOrDZGDvhIWhaGFd80HMjEQe4iY/6LPSOt0FH0pWR
PRe2KqeW7Mg4RoBSGgVC8L30DnITPYqk3oO0YKAEyic3WuZhtmmpwaaAMKNLsARQ
nNn/LTr9mKBu4/u2/px/P/zFFhCuMtIhEG7KBu+D4BnYSv5zQNnfbJPejLBmXm1o
e2KvzjddwMDwUVfqqY5aSf1oIXakrXp/DDmUQDKoYe6huDUH2sdUZy7oxi+q4hJa
wJndSAenPRjMwUcBt0j8ext+zMhXPSO303CmMGp6FcfZCd9ViQnobcW+fJWLmn6M
3R6vYproW7caYvtHQaOBig==
//pragma protect end_key_block
//pragma protect digest_block
aFgjWUO+nOLqDKSmBFkS7EuSUWg=
//pragma protect end_digest_block
//pragma protect data_block
wyquIFLtgDR7/D/h3R3cdEI2aOcpRlLMAd7HtByIFI4rme4jhPqwGDY9/KppTJ13
mpIXpBMnzsLDYz/fz+98zVhGe/Ej3LWphQ1lFfDBl80Ah5ZJ36i/lonjIp9q7BvE
cAu+tX78NbhDRvTuT4/Kn2nQspdpspv7fZJAKv8CVmbpT+B1uqObROFe49q6BUGq
s3C8+8uC77ohTyZKTrKqLxcSOrXVQqencWPN4F70nLZtgWK/N1SlDQba041TPfQ2
8sB669TWio01zvU1whe+A+ztQab/Q0wHcNZF+efSjooJ2f2OJ/7OAz6WQyUqMTFo
e4tfbXWujVjA41wMBK2GlpEOoV9qskoOuvLg5kvHkfz64pPAFvnPDDibnuMk3T+T
rI7kT7P3rCy/iA9+QSZMuYhx30AmdWGmPB9uQMYOwho=
//pragma protect end_data_block
//pragma protect digest_block
IbrwFRDp2fgjDPVzwKUYvm5iQpc=
//pragma protect end_digest_block
//pragma protect end_protected
    `include "SS_SYN.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Ai4KYy0m8J2ZIV6wpVyUwe+V0TdA9gCNZvw62OXky5HLJ4X/LHHbtXFWrygiJnnY
NdxwH85aJFWZhEp2c8/lBfs6T2Hzf1m9aAGlBDyPhCYUo4+d2kf6cPCnQYqEsZJn
R6BqUf7XCdMfPXcTqvzwl2nz4Loyx0FUY41+FnItUAS8SLqEWhPxpnQZtCgXZTqx
eEeecaitDscKjWmYwuHKWcX6WjPrGaUnad62LWULKg0jQIROA8KfczDfcsqHqZk4
HCAH8k5Z7Hn95p1ZgEeVmprWQw4O4/5RGpdGAyeZJvx9Cw5HOv8wBxPIi9b1TUQy
RGY6MIwzZkH2eLufcpuaWA==
//pragma protect end_key_block
//pragma protect digest_block
frlDk+UcdjP9I9m8CciYU44d2gA=
//pragma protect end_digest_block
//pragma protect data_block
D/SwM8vOUqk61KMbbhhp7dFFbqYhIWBQbPG6hRHbLGSPJcq7sR+YzCYsss3lsNxa
4BDCWK34Pu8KxWDXSwa0YK7/12dOH0DP6pdeuD5nlms0XbFFpK8po/UpEU5Ngx7z
Asvqw4PPzOhtd1hu9tIFh/kyuHJnQNYZtr5y5RUEes6b/PBTVEK+M85fq28ufCWA
4cbOAMy6lkxyLqJwFsYznFxhu3tlJRGrc9JaJwBOovJEGvojBB2hV6KYUjd0rsY8
l6p/PEzbHs9oZkb6tnrQpskeua64QsOwe1HTrxHkHhdoesjZ0jc2hGKTIEAtvY7F
LNarlU4m3FiUWgg1VROVifmfeYkBFR11xs0avSlXHG3GnKoBMn6h7NAKdyZcUQyj
53cR/Scp1Owr56Ac2qTGbfVwAbjQbw0yNuIMKw40LwTrYu8sRw0VhhIzWo+en4mY
woWaCaRbneLtC3GOG7r6cy2ceBzaqknfrXaALdvZgB/d1k8iyJzURifQDOV8nDdb
mUxyU0+/L0eZWTr+ELcc2CB8NQtJ509+1svSF4wSBGT49uHjoDfEASX65JAvt/Ju
0c10LQ0H9pp5yc5hnnu0ZNtdcXmGagCf+9EhUrKovrCTjziCMfm9SNTU/Awt511l
Z6HWfjh8/hN/4UP9JxJHgtCLgOodtkYxJqWXZHZfg0LtvIvA5zsABOL7XOQdM3+S
uYcImEdcPQaAfqlWfjTfvfDtDudbCcOvOHxRNWnak1L1x7/DPHFlV1RJO5O60Xi3
3rpt9eJGGnhgNZwmuTEJx8moth6UKj1dbSjEtcc2cIPlGMkgfuWAHhlM4iN0fPfj
7pm/AydZkQ61eed5JSBNB2iav8mDtClMpmua5Llwzz7+DIM9M3aX/juu6ciow078
F4vPs2zoqC5hcixF74FTB9ikum8QEIAzNhiY381rD0A7sxbPk7TeqqMydCBesdFo
jpk+AW+ss466+UtfTYU0B8f8szjtXnNMyeScPBo6fzlc1k7ue8AQc4Jvf38q21DU
9cTrxtxgPx6FHUujZOCHr5I+FY45vK673h0pIHDmaSquPRIPGCHNg+T8TpLWyvSH
hs5/ZbHMu14arZBhVhJ0W6U3eGu94T+jIh4464OO2tXgjjEburN5SXbID2mCNUpt
q2CL5v0DAUkWqQJn89XrOFx88zjgKbTBB1jW1hRFmboTswf4ze6dg26rzkICcr4v
pWuf/u1MKfYebI7yJD/Yph2CUgWDmELAD3MDjNKraNkyME9phTXLm0MZuvtDtwHl
mCtdXynBWtlcQm7q+pcTL8f+ebBu3mNX/uo9O4sBTPCSHgi8Yo3u+TCoWesdHrxQ
Hmerorw0zTpPfiMUQBHhaCG/QYZxLaTciDTN0I0VN3VpCIyL5i45EhoV/ayz+T0X
9lpaxUP3g7Q3nsdZcBm+P19fspXqTSgJEvI8kne2x8MgaCIB5PPIUF/ywhwlTVvG
g8PRMyq7i51brd4mOItwxPbGY/QsGIVTyIJqu3S1ygh1jcPJhbgx7V4lrGtpfiso
Hi8pss82yk0Fz+u0baQ5nkYtRVsT7ZrcRDqadm8wUcS/fqkJsn3cnj7SygnqOJxg
e/EbKmGq1TgRGcy3q6axvLzSOMVbyKRAjPlyjFPcYbr+AQhvo0JZnIIx4pQPqcYQ
pIuZ2KvmR14LuO3Oi8agUkDnPSTceqgCh8sJdrEbFup1pzNbK/RRXKsgxcTZy+t1
7WaxlyeAgD6pZ1ku2+qatbRmWasfuv9oazsZaKF0KgW3/rxPQIXKjP1YoNVPSH/4
pJjcifqZARdAiin3eR4qzkuyVQrvkLJf66LISLyS7lwlKMIbHPiaqze/yWlxSNDl
gsLhMID4aBQzYQEOxxX4vBQREZyQ8fUmfp03I3itXYOQlQJ1bS3HAZ0JVGoYM7uZ
l6dbOvKyZTfCmci4a24t2CNJ8yfTvQksPWwRtoM7zAiYcv7PcqtFTr4PydjhZSZt
BER0UzonHmNH+ddelsc1ZG2PLUZ9cEJ2FHf43lIKcJdF3RwylK2gZcnFcI9aY2aq
64x/u1e42NJMhOq6csrsH2yH1628UkOp4JxZL3EAiRLwtvXNTSKqE4y7PkDvNpBr
mjSKWDACqK9Ap7uBWawPBTfQiNv2rPg95rjdpJQYaCmkz9wZI4erVeRG6/F6uLgs
cS2AS1NFv9C/8AiKvUpsJGIR/YhfYuF6lxZlX161v73G/bN7rpk7u/LGOxAsV+t6
CzgiDsVFQbzSKzhh+9jTPJGFPvpLe/mxIEKC7DalbzXHf5oBzkCyw4rJHxGJnxsr
oy7aAnjeDL6uvSnsBkOQAABIIcwC1Ofp4ZxBr8apOteR9n2Uq0sEmnonQzDCtrBU
j58iV+iUJU5UkwdQhISFjUWtHwOJbyScyiIN2Mw6Z65HA9OnDVaRdvgLGhzD6Wok
iEJ8FZuqfwnwY6/WjewsWk+HgfzzGcDxNziAhtiYc5gC17u0m9NIdeCC0U++5fxJ
2bsAuWRgFmQ0t9zKEDr5SVilOaWHDkEklYGfPXwq0D258B0gZY/26WdunXnSH5L4
49ddAEXNWRKzu23VVJmyXhmqi3dsapiJfDJ/+jmkJXe3llavQKOKpgnr9it8QP00
KAczar27vcvMBhC2CWsaNJlYncdDDHCvQ+HtW/YqTM5JZaApS4N+6P3puFgkHjVK
c9HT67RYV0hAnFuj5vwG7XTiH6dNXhEP7UxK8HA+Qp2HSK9xAMgl/FXF6SHYPZ1d
UihXkvv5BYvBIpdlfP51NsY1I3Qz+phs/7xyvewSLDPOWosAqPyrMgiyS4p3IV/X
1JczChKg+K/q3dLlKfqfdwaYfXXFjwIODGrvV8WoMLQy3XXc3fl7oNkiPVStBQlD
yNAphNaTXDKn2AJpR5BQS+QGnerlUHQIwFifdgoL9n5SGeplf3Kt+2kx+jtFAqWh
G0bZPOYTMwacDOaOvk4q4qRBNOF3VY/o9WBMBxAx1egqfpn+J+GM404c7xUK+c2S
cQ6p5TvkusDhzH8gwbDH/4fcSNp5NFEXTHPH57HCE46x0lCLfnyhJryoEI+2m5w0
9p8P01wyZFWe+3qCtomz4AtrIfj1BILof1ibnAfQZTifOss3SIMdJQdoqrpC+KPQ
E1XMU3lScEOBfT3cj42jRgD53Y7KPNDu4gBkotuwWEPYjopEmIITylVrRUUP408r
aQxZNB4DZBYLJaBW1Au9Ji1dS4paF+Qf5D6spQmiH1KsZmgTuGhXOm8qtclVbh49
nUbH01MGQrZF6leKE3PVwlDX4qXZId5jI5o4gHpO2YKgVMXhfRaOUS1W5Soo3vb0
GwKFvomcQ4brLSB4t3OIe7MOghRNrcyNNHoOdYICCBX6kRpWx+P4eKyeFwgrxi9r
lMK0ACJ48/FjSgCT+NuRZeuYcErKb9NpEktDd9X06rF5DDMPKbIaxU7Jy6DWu3mP
0kqJiUC9pI1LnUNJco41vLN1LuWCz2u+uPcrK5VKNgE0PlhjwfsfECfJ0WGi5tGc
Pr/12DAugfe8PwmYVzvRp9yZ6lTCB/sp3vua7EaqzlDX4K7j0cjaGTnIaYRWZW2+
/ao3EUnfjeEiqNbS1WHZOPuEmQ1b/tq84Ab1C1cZiYVHNmUQ3+EVBH1JLEl7HsD6
k3ylOiTDxoSPhqOrpfmWcB2QMHGsqJKLgKjQ0ky75ubdM2keb/pFgnN1lpRHdHoZ
YisPP15UF/RRBtIee3F0Mr66hBqdrJpIAZhsv+DKjZAcDjk7KuYev5mPaO8ajbk6
ZH2vpKSzt/ngfzEGQWYrkrXaYkneYyy9x+XMbLT5qhP9d+Mh8qAgGBWNHDwEu5oo
vQsuuCDOwOXubwqlDQ01lPxECdeXzen7pnX6vwAPcIypohawtd/VXoW8rHu/LOhu
Ue4dv2luwriAd686sLgLqwmQXWSlrB/hV9yB1GoDlr7nVwk3hrvlg5OKI5PEARX0
0J1oFF5VjZ1WgD4BkjYD86l9PWfk8eTTkSLmxRCH9FveGR/1iL/kH4zUaAZnIN34
G71w2W2vDlgdseGMXHN+wUlQxXL7fGJheauRKkGoulkDtqAj3zTzAqkCPqH98Nzs
6aOJEPM4y/r3S0tRhtLA+Wrl+D1Q8AmZVkoe3+DwNRXEco4PBIQU4KJwmqouUMsw
SrJX4ScVbJIkA8DPD4zUNoF9GBeNmQWzu6GeV3gVrORiw1QPSwe/bje62wo91+J9
YLiwrGDzUAEBB4fXgI83apMHlW0N+UafoeQN5xRV5q7TBB/sfq3w+VhL8g1Kh+xm
mmo9Bk3PfcJsBvUGKkz44UmcenQt9DLzw1SB/zgPgcQisbcqaIZDkosq9X8N40JP
DE/7P32kTJnPW7fy/Jk4Wa8CxKEoag7JPQJI4YUF3TW2MaRSiKxsyTqKn37fpANv
JOrzblelL2p/O8MOUcQafe44vQZSKzD9DS2VSb2y0TyVru5Uz33YsEoIUwr0nnEt
BqHC0zyHToN0YPDq/g/T4vKTyfaXbYMpOtoBu7Ykz6ZXdW11eazAhf4WK7WpDVtY
A/f1rVbnO9qOYZKYqmYss0YBwzat1TGqJNF9j2aHhRPBXo850quznt9XhE5UG1ja
bl4hhWZmaT5hWE8lOOypMdk/YpXMG8pqd1fUxDylCvtumrxogNgbEIcFXn1ejAUx
EyHKfkRMyB8zYihxocmgUPzkYE7Be+AcWOJ9mwz2xoJAwdvFOuqwBvFg34z2ZsJD
cZa1gWrxuKTvyNA6OgJy34da/J8JMuquXEF4PxuqEuke/Fsm77F1beyywnPq3x/9
UmAUg9/aG39fct4wUQO0N7DWptAFlux0HLai8MIkOtBMQJvpkDTTIxLKycntClsa
ziIqFjTkUi5ZPZPCbAPX5bLMCFNPNMsYn4xXgFepV5B+WFzgQuA/Jcvaqy342+au
Qr6OcyHVBQHkuVChq6O6kSstvFnJ8OWKAkcbkAf50hx0L1Yb+AKhPm8L0g1Tmv7H
sCKaIk/5a2NITuX5jrVsaiAXZEVYE3rbFmS+VnozyOE9iRLtZ5yK8YwnzH0iRKfp
lspcNNnybE0lbSQBs1flEKS/HiHOSy1T3W07p8O3DOVQ5KDYXKEQxUyTo0N3Nykj
Ph0B45hNHab7YGXBbRtmcggeT92WOBcPZ34D6QY3yvSbVbWkRjWOcrYr62DKlpC8
CFAiBCNVtYWharnvhBYFw0YLTc+cwOpF6T3a6Gvn5VaWYTlqQVzH44d9v1WaR3G1
Maszww3wZOFGGeh5TqxvDp+71JQsGNag7AVruWl3ssvnmxc/tBaw+fz3MzrZAf1j
SDMyi/GZRmSUV8RibpjnlcQhqeaklQeBgGjgKn9UZJvRCDpOD2r/HguY9x5dtnZa
ZGYqdIJ9B07Btj/AwGoFvPPoK9KbI1xe5jJBhaxEkb8MnwGgKcCQxDI61ewZc41F
kCYFVqJpgPVHysMbqOVRRbeF0cfR/ugkLcFKXCeo7PPfnGTTroN5d6kyuGfI+ccE
OfNlxTsLC1+kDCEpuI2vnRb5E9uINIFIT7YDp8LbQ7FrOnR50h+pwIUawzesgGbr
kHSqJBviIlBGy6oQFf57CvcBxDeAPmg3lo7LOQ4qqtBK6+SpUjZ0SRs/pGAM5X1P
jHPxDOyhvLJn+XFIvaY5TrwOmNIuuXFANJGifcIMgi/nYVurEz/AafjHAKjHMat2
QK+7N/MIUv/9zY8ubbdFPVUttVYPIv9LnPFbWtICC6etucgRBpu4lzHhMLV2Uwg6
qWCrZMyLLviwJgJMUJQJPLz8cF83n0L1Fs9qXd0Lp8Blq9e3Sok/p1xn+h7PsgT7
RHiM/OxY7qDnCUpMYNoumAUq5midjmwzxTM9tAEHISr9HETNgIGwkwZJQEtIh1CL
xP+jiywaHF5jB9iEfnnOgZq0L4KINRalpaGG9L4XNfPswkchovrQsc2Ri9IHJ3Xl
10dyBAGp9HiA7Uw9P4TEHO1QSgIamhXeJdKdXcuuPI2xLQv5ZmS/qfQgTiQXg7Bh
LeH4+W6Puja14zx/V3xLx4/l5kiz+JD9UPAfmTW+afE2JvOoMrPhqzIem5tBfKSn
bfrg8weL47YUA9UL/9dIlH6kfXcmfyz4hfmoLkCYBM1LQGHFySrAU/RPDEs6DSlp
pknwzDGy6ut13rRnoNNO7pIzaX3WcxpADNuxAIvQvvGo8+oNoz7IFMf93GoW2qWQ
0CnamHLmFm4HcfXQ0Xt6RoaHcm0Qx6Ef+2TsXrB4gnKAxjMlWRDgK7qyRMtgwgGk
qyn/jVSn/rZRv5mJdUoOaQB1ESNg/F6P31yC+SnnLPeoZ7ny9P1CqEXb0uy49KTg
SN94QxDKNC2SE5es8DvvdPik60UMqeYZSgbbVPA/R9V1DK+cH0JMOahBwBm4P00c
CZRWbVLfjV/sP6CAJCz/0GJYTA5V0zvwSYVmv4Clo7PsZpgrWXsdeKUfbXFhKtnK
HzlcQyireuc+9xWzF9rJrrKSUzLEkqIHMlj7ktRiBH0aoBSMabD1WBggWsDYSuLa
Bj7QG5ejZ8Tb5K5Tdf1AvOAxP//o2Cj8rJaXBUhU1df9pLtFrL2B3biUQ8VtYfev
ajxGN9kb0+M3W1oKaQnoyjikR9dZ9nqBLsZ52HKk7sgdKff04AmmwlqX5vp+liOP
hBHjFsbq25IMcC782299gGHtZPYv0XTFpffsUWba2j+FL6zx4GdL7JK92fYA2F8p
N15oiLYT2uT4GCarJGoQh2n4K3QNZNaAGbf2o6eV79fUrQI8cuzhm7Ac3L3/EtF4
f2HvwBfmnjVN1QCwBj1k7uq/N9ospsTGDKs+63wiX/vUqS0H/ihdY+Ay9tuyALjJ
oTv6ZNmAESOFOuHXkcWIdCPJWWxWqzFP+PET9uNXJyq3MIZ1fUk+116iLDXCExgP
BjPvaOI6Hc6lpmXCUh0ROPICtx9sJhPxiO39IH91xLR06+KmG7lim3P0DzTlUQsL
AefyotoFvKXG63VNWkw9IG0asO5b90Exz4C53mtfuG0K1S/KDTRLH0f7q04QiMvn
s5dxzN78WqD4WCSFh8p/NZDYY6N7UHTxCp+u3m8xS9umKTyX2WqTHZyv2q16r468
fMcIs4J7BhwW2TmmwM+zsdCiFbjiHBDTFIBEW1pgx8RySPF7TH6otoZxRDYoYqSi
Cm5GA99vVACewMNt5YKOsqOUIuJUT9aqtXFJ60SKdaIhVN2K4zbjdZgnM9ADgobN
jofgkRjqBhgRVHf6HfwQCzfpnbaJLZeE9vx80tCgoiVtg3DC9g97o/QOwwB/n6An
CMdWk3wPB5KqZa4Fiad5kUTMgJU8k/27zcSEuZaxpMzoS3/OzSoHie7v+PNQ5q9/
5tfG5SF9mc4Gfhi28ClJPARJ1Hjo+YWnqKtGcxGky+tFI/3Rl7sCSNysiAxOuBIj
1mWUZ6p/gsYYjBupFpj1gz6ImLjKVg/2DI9u19VHnIwuhqEtuKaCgmnIP5ind+nQ
lL9mvr37VYqxV0MDU/SGyYcOvDoRxPe2LoK6N41TNBvBLM/F0OzQQJWztRqz3zBG
H4cPy66Gb/xZ55KLUV0/TRAt9VR4rjnLihC3uv6OCO83JfN22wQ9j7nBJ8mJnxc5
eBynSLhk+i4cYH+HOBJkBpdU+9hg5o5i/tDgm98DB97WeGsFlJrsIYVKFnx8Jivr
guN8uX0n/HI/rTUflqnojSP/y9pfk4fonKH5iGQPF1qMn3+XvJUDQSWS5ZYfwCfQ
lQIALAcXMuzFVbRfFGjY+4tj9TUGRDomsUvWOJ7dOL2ExLfZ4YzcGdp9D71qMDwR
KKgX8XsSNo2ydw6uaD2VVQQIKibhyrRJ+Wy7Ff1zN94rAkIS3SWRqUh4M6E4rT25
bp3bGOLId9QcwnlrDem99uOmj/wlR4OUrwfZQX+jgJwUkbIkcaSrIPp/JDjtw9vY
lBI1sCTbI6MKVHCErLYVcFl5B8yR5aV9507Ah/4LM4QYmk12iHOnJq7CEAKGf1dm
AqFFUeaehjVCKr4Llor6TGUSv5rwwDBVDq76hu5QjJn/5ueQaPtutZ04LJwagtY6
Fa69+SEWGOdmZeURyjJkluIl3ZUjQ5zU6B89nKKvUJwn76X5PsuQC9xVJ13jqef1
dMLPD0QuXtOWOPzH7d6SAB48CSVQilx6kdnMSUzQLNgzpEPbzCP9nhu5/xMPrlhX
Tb/+4IsZc93b/HjLko+KPwHgh6sK0EOsnx2oQx1ebRJGsNtsTuo2Ip5oySMNAfF2
UsWWXJliqwi7huwsqIdQzZZ8p8q9/zj8ce1MPLi57jCKKtqlvBu+7vA2oLhB8Wyt
cH2ICi53Q5Qo+KObQXxaQ1K+bfPagsERaYwzKpzRNYSf62rHwKeftFdIa67HoTaD
DV1mzAwxfYCI/aPr7dazaX80AHwGLG2gqDtw3qfbRhh7d5a9uYYkCazkNVU3Svbz
CntfnZ/foivIflrAbVDGCX91ghT1T7qFySy5twIfVLC6ogtxeVjkbje3mG0Tkno3
7pBymvYRJGU2GxRk6FPKgf++zQmzVYMPvUPXnBKXfBbdVibBcgPpsa84lDITlDAW
WVIqizjk0WwR6fhTPDp+Od5dzTawUYJMHq3TD1yf0nG4kmnERcUOzq/ZhcUbVluk
Nad7T2Ic1y3hr33S6bFM+pVUQNHsLVvzWOAcuDV9fQUZWmDjqNgc4hQAX/MkxnmE
CsXVl2tR9fMz1+2/IgOVuI2IjI3IpqkRImuKWz1JKtwDS0M89vyl8UPDGstN5+eF
sXjEaQE7vcrQIaYgP+mGasRYVQIoLUhMTjmeaNpL0FoXZ4CxvEjFKB3GKk3WTl0D
58Ik/e7EV99CWvH5iYG1XkDxQFIle6iJ6nAvcFhg8bXQLo0IJb0chZY9Zv8U3u1n
FfIc5TOLmeiExVS/QKakGKuqb7gNRzPAHK7IbUNY26As2QoUCQ0Aapoz1hGPnwQH
vPO+D7W+S33t9liFYVi0cRp+tnt52B4oBnsA8XVoa2gDbyyvTUH2/mepHtRiSpHb
JCArovjDepOzO0UJzi8hM15/Wu1dcsc3QtUVxGdRlN8FSN9kE2vksvCnnZcXpwVf
HnTlR0mfIjepEYyQoQNCW2qnBNxGaOvr0OMfDXgDb0zjDi15BO55T9aXR5fLRfqV
s5GLypxSwGmmw1oj/D3Z6ykcpeWGBQN9bxdUXU1BMxQ7iyp4DtXiGd5FYfXHwYeA
iwcBnPoPVDwTUHh1H4NIKuv28HFiE2M4Tr2gHCnxoL5wx4sSN9mppNXuHMPVX+m7
0XWXrEJhUMmvkSf7cawcx0xHAvhiLNG4jmY6w/axf+MCTtGrVy/PQBRKvXtkHL2q
TBe0rVL3v6sjCbUq+ngYiTyo5Za2rykargigi89dOdj45c9ZKh6gA/p0tYXK95tZ
l1u5TSkZV8YVISzTz4dF+qBXzGM5tUiqSFgJ/xF3tefHwkdDc31cZhZZJzYFLLRh
zS7jS3IjrfcogCE5oKGI6K2MFdbwtk+YjOR1JK9QbWBdCwZRNfUV5ZDNiM9YIt7O
ranBkh+GAZ7IYRLiaAc9bwg7kf6pNZ1MvAu24RXPbkIGZ+fJUZDAXHM5zCdLjCtH
Od0484l96SBsDLe7Qt6Jjs228m2sfij6zFTuV11H4wE7eHJmB4cHVrCY3kjLIgu7
LfdmIQ4VdzIuI3tQn9VRrHWmM6GPNAXhU2uX8rbvctQlnNMsYeO8hVdcwPZ7obCg
c+C1aIRwUi6GwfPil8WnszrjFNFrstBmVO3ml3ajDIH7NM3JK64XY6Gto0P/b6xT
djuXggoHiRVOubqD/TQ8pvAIQivyxCm+YqYCl+LmagUXOiJDt3cumluKJVlyv5Sh
l5OP6XtHAuQ04A1hZ+I5hGA6LqeKhHoDbBETh0OOe+ltD23+sUFKnbBcdJtDms+I
AvIjd3pP9Yt8Lzzvq+p2p8AFylcuhg7D3NZDbAoU8/xZAwbP4PsqM2XuPfFNrfUC
nEh6tEP2zpiDhMcW3u6HUinOm/Bt0oiZRWW43nAgQnqZR7V2vrEqYpKjXweLJoSK
gtMf+Ei/SqPztwj6uiSIlsQUWXpNd5IGaZWjpCFptsi/O3bwQfxEjoGU3hhJ2oZx
yEOgNCOytzRsy0RmC7WMeSxPIDtoSwIbw2Ynf7+xZHil/614pwBzfuYZ4SH9eTJx
9esqXQvhFebWUwy22tkup2rjbEj+Z8Vja8WqQW5bzft0NueljLARNZUqa/3r4PaL
JJboKBD5ng0z7gQx1edB/yfK1/OvXCsJsSgHu4JKLeorE260oYL0yd6Pi+mGRqGQ
bXZj8rQpmhUii227I5kcUtAu9/Bu3f8npC1XBfeuCu8Zx9WmrYuCvxXgJ9i/mMTg
Vv5mT0a8NQRUpVvDSwcIBfdQ+Wc2el/bgcJDpOFKqxERzaSaNvLna9ExT34Lfjup
Uaf4YnE7dPv2x7VMg+0K0ulgUqjj1M13fEEb9CI1CXB78lwnHJgc3cbFgP44vr6l
hyE8fe64+RqoeEzZG/rLoHYic02rtRJgaxO8BX2C2PXDp9YGpZKnW3CirmTSAe49
ENfZ4k2ZkiSMv3ju+bzdZPQZwXPyV0QEiE0IOfOQ8hz6mElHGjpgKbWtVYx5/Jdq
/pZBfsrNqep9Pdk5sthZSbSv4aKfDCt5QMhceQpmADlOlEmdTCAeq8Wq4bDT8AO+
Ci8RghDdYVE0zNWyRmysK/ipJrp3uk2mWRizFfuvt8d16NCRuozL1wBU1bbqJ3Lo
bhRIhD3DgnWaupiCajcoxGVhctE1MfPLUedf2TWxVs8e4JGS7WcSXOMvI28Plygk
IG+SlV73qS4OEEo2UwKse+FM6XIvOqzIkLuvlvpqQzQrnlxySpcsTV7Z5lHOF+/8
YSbJtHiFFPZJ2L/yBKaaCT4dl2fL45OuMKZQfZh1aZGKtIplHOtn+nMnpLz6Uxaf
4TOUHWIFJDYXN++5LY8gDY2PwIAsaRa+2dR4ZLKkDHe+LLvLnfobONu6L61EbMVu
R7+wU/X7k67wiksx+J1DZmvCjk8b9LUzEaWA/ggfNWZf6KZVRMgAqwkUcPTMCt+1
vH/3RL9P5HzbOVUkNagCs5abkvSxwa0sKFQJnfo168ZQw0QsxjLZ2MgauQXt4Vug
wIUwsotDc8sIOJLfK7PMZe/BWiLLzOo0+DMUAJlEjAPUi0hQnplk2N4+189EM0F1
w0H3ta9NoNeppAWg4iaYw1UUjFa0lGo3aBlPggJFr1E=
//pragma protect end_data_block
//pragma protect digest_block
MpDqwNjKZhrMYSfc5vtFjyGFy5M=
//pragma protect end_digest_block
//pragma protect end_protected
