//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
daf7axs94+08cQKOhqzTej9/HIxIIocPWxcVW6gNocZ0sVGZZTWED+SLUkMDZLTv
ktLZD8RRxiTSOSG0socc8pCsuyQbO8o19jo50ptth8GTEKQmx1zEwr8qHnDcydT/
wtcOutjUgAFU4aGkD+TkvHeJoa3fZiW03cTZ9WOgW7RN420CU4Jqpg==
//pragma protect end_key_block
//pragma protect digest_block
TWMNIr2ED6SpPChwrzRL8P9yihU=
//pragma protect end_digest_block
//pragma protect data_block
2Zz1rMYK4n969bWxPlunuYtFrLWWJWK5YkLuI4IG1wzoCpro9IGg0J4udfMQUB5c
n+xn7poo7g01W7DR+QQMuKuLtlOJPWH8t5HplPAQzOTEqIWkXQ7uCX4yy7FtX3wY
Bid62GVM2Ieee5Cikse/Sx9eIC0AsVyZwJybAJnbUFfIjcSg+zuelKaptw2uf20N
ClkKX8SNLBfhpeOM2VE9NzGZyhoS1oD4KUw31FQceZxZn7m116/TDmULNhcGFjyg
jR+BgT1CuYGnxt0Jl8cnYV1AV3l/tav8mG1ByCqmMIwPxww0hvj7ATC0wBX/ut+Z
zTmJeLhtNlmAE7HfUNKcfVHFNGKMpMdrl8dAVz4mBKWsrNM3W0lo8ZeNDBG0aqKq
AGT+gaPKT8XGraV8mgEpTm+ZaIvAv99md2uNGMPM57hds20cmwz1mXDfjmCSLGt6
T+cLYsi+cX3eaIZwRvpMu3DUs6WUmmYwW53j28XGgcNaf9mBnJhUnLXv3pZvBMgw
dspBKWLoPqNc7e9ZiP6M+Qv/nO9MEclDkwlJKmW3MD5OS3lI0DJjknvSopCPbQNe
DrZ7yBhHUrOCO63eIraThfqYrdy8QhNNjiYicaQBdTwiVbE51kZw2ND3RGwg3aCs
Lq6A/lLrcOobSezNrg/XP6VBbXSKWR8y9k0IuY075uioDz9piIfOGkFVprkkB8ue
YP1Er5L2hyMQdcx5BViXdU/m6gp8+CODHjGuUDD8AXUga8RAJp8Dy4o4fmV+e2RI
PL00kycPvAVxGKcEYeF9o7ZvxFpXDdRo/XLdGMek93OExLUY8CLXfGunu2VtG6hG
xo2LGFyg5UFJSvyyUn+oPYLU/Eb0MxCxnzbWzqPd8N2spcUCxRnJbX5OOdPyP8rN
gTelKbMmm/fHcFkjYL8Oz9r+6/cu6l9ZtXrbIdATBfC9NcLRjfRtIHalfWJS08d1
R8dcm89drMWpgAc8J2VtPfjOCJVRh5tjgBJqds3CX2ox9Y25z6eLTrC4hQWh/ym/
V4ef/Pw3t59+f9MZmqjUTXsDsGQ3wLck3PlyTsr128NtvEFoECK3Dr/MQLhURUU2
2erbsrTDpKKonlNt0W2MkjkJFB9KOqfzJWkeueELppX9ejFMTOkY9oI/GnuuWhKw
Dyytc5X1Qj+CSzo7VN6492baXf0OlbugesE8+/M7F4bF/NuqjGfV6fZdHVf01ySj
GBrj3sAtXyFQDRsyYZFvcchItz8JMSzapCHk/zH24X+KHuwruipyjgd/JlG1TZMQ
pyVASLJcCyIoFNGgfZNchzEBQKROqp0WQgLQm2h5et23Rc6Q63gmdnIdaiFJjfpq
zzVfF/RkvO0kcUwN6ImZi61hFbSTmpJUo3rZD5vR1CaHYkpmwI/CGPKM3uxuyIyE
/YL0EPhK8Z9SVphRvPFtNeVwTKagtZVxTr0Tdoo9ZBzdUZ8dGnOT0qtuRJVk4eNo
T3c8IS1JWjXAUypFsuwFJB9DVJ6uGEIRFctlRo7J0xhgSCExVhxyP9EkOS06NgR1
ZM9TtuknlvJ0hpM8+gZHoQblHKeyAKKPdjebXD7pO7WvHmJiCTB66PER7apyrD+1
KNmd/VE8mYx857lIU1q1WHuL+JYbQsPsEr3cDSpTMnvfKlG1Y2z3MweesJueGFdz
DJDFWtoy7lTO5UnGPQGPzuVj+HCL/LVunvc2nSEtF4F2B/9oCen6g9TrxvCP19Hk
JJGRr3NcmehmPwmQu4cNG2ShvsFrzpCWdmtDHqVTZ/WEaae8pIG3rSwfkgffqBl0
lw993zJ9u84xoxzilAp96XLChIKagLfZVawU404fZM4Sy+0oDJlGSEM4G63GAha4
ULv0w/Mjc5maH/uqbeuRXfBa8O8y1BaL2yN39+Eg2afh/jQ4L1aWYae+bVUFUreq
5f+Fkwoy7nA2oLPmCv3YmYL6VwmsgRFrQT0byMoQIthTOfJEf/NvIkqHyevz4qKm
+M14RFBk3rKCl/ewsVEqWae6n1Mv947cKethXyyMCqdS/Xn2Eu2rZI21a9iEyXzt
LeUup89OK2uhP3OaFT+9qxOZ3N8hhUzokvAhwxZbbmthExOdjLRFhyQdmJC0Yky1
09zHkm/UeHOKOyAR7oI+0WGGtnH0EgIP05Yl8FoVkuXWH4VSmtw8688TqSxVg7ga
KUb/Jmy5fBwHSM2y/xYoLZ8/cQjqEe/wOmAgn4u5b6kIIaOejKvpOl2j4gMB7Teq
AnK62ZgPvhonZRtcxUE9X1uI2Gvc4bEZrFpeyo10xgIOqZOd1yDG8D6bZuzcS6Xo
teXu0vteKr0hNFUAeHiKOaKQC//K5lpnkHEkbBSco/XrknMx6XNrUpalFMyiyokC
hUUmnTL1U6Ads3Yh/3Mr3fVn1Zi2gAtvDxTOumJZx2M+cW/Xr4s3d2v8CKk9/B3/
uof0KBbaYHuLEg1v9M/yVPVXSmkYYz/OMPRV4MVrKBTolXsb10S2yS1pRLwUs54n
pcbm/g4lF1e50O4vzH8dHWkMWiQ9d5C25oFulck3qEZfRtMfizPOM07zV7K1g38s
Cgr6EvP7khQ2ZfK690D+8NUjWuuR8kzt0O07T8r0cxLsdcFprerwC55DNUIsU18+
3elOOojdJxqHRxlQh+OP/kiAMFj8j1ddE1+7ta9BbFmxkcPb7wbNVwUGfsbLY9az
IoWr2/Tez3C3dWkwqEjIbEo3da6Z7RdDGdFbm86lc7tzlfW3BY/5/aJgpMZTaemo
Pexo5iQrc8K/NI+P5k659n2W3rUd02PoUSaOsOPvisZKiQnLz12TAAsD0xc29xP/
6/BSL98BQZv6qLVvQyiu4PdrdLOQp1i5oUqVviK3yB6+Jya+4fXigxzBbuHyjHiz
LOQrhOh2wwUuXCZX3hoVhJ+G6xmgO++CixYGplGF54VzjXGpRAn5/9+851FVTrjM
cqXgj7QAPmszBO0wxrpMEcZQbvlVk50CNexCepPRxG5kOBzuM7t4svRc2fPT3R1z
IjR15z42dzLC7PX+YnZzmpzq2aVwmg4iaF0lZYMtYA2ugTNsIRXZakAbGNuJXg4S
TtRV9MAxMAYrz6RqtpRB/wCu5+LmHyg60WlusP+VC7YzeG9oNWkOJmDhUdnX8sOu
WBVUvdqAzko+6ApgG+V9wM2p/175xFOhnA5UsIMMAvNioukTMBUvqWDGV48kJOUv
LGrE57rq/dW6AQbZGfJJjrwMkIippwdJ0uscnjtoyRhBnGBj5ZZB0wbHA7qY0Mwg
IvoqpOMcIFmA2U07BpjU+Ej2+CJDLf68Lf8zU2UCLeAuqq+0Wnf06TylUinO3/+n
Edkrvftoi0LsJITtVef4QXiHmKd9k3mvT9XsjARFCf1v1z9Fq3dHdj+bDFslCl1t
HqU9WVhIjvRUTlnuJHDL4RQuwLjti8Cmw1V7b8Iru7Sb4n4gysDfZySGH3H28rmb
gu7oW9VAv4qQigbLX4SlBbMeJ5x51du9OkbPRfrFm5eSkd1tH3+rjhbMmDc2eQCN
gG6BCaF9qo4TcSvSkETyt+xDqv+kDxM0hiaSV2JYjJC5TW6oO5NrZdZdQneTYMgW
FAwHoc0yqyMBsDV/E3b5REqCvVxFdH1ZXGH9TVJZ1Gpoi725YOwa+Xz4+YaOUh2M
Y3iiIzunOlth1g7mOoliOpEn9e556OD+DE5oW5FQ51NveDvh30sxVtPUr9XcOl+5
04MyvPmju7ho00ABabT4/7d6VcLycmhdk3QQiXsIkUYJ7q7d7be+Yk5mMV1/pIRV
YpVdOxtaWs1ftJ1QE57YtxiB3UbzqLrNWnbdNI4OTpusG+xrLI3CY86ZvcZ4S6Ty
IxqvtaSwrPhiHqSkCKyd1pk88q015yT/HRBcnRE5/BHTLTB0E9X0iuwboSDpe9uV
cnLIR9jSXlXN03d734BX1FJ1Skeuvbvv66v8uhaUm/xoEJyIvDC78KuD5q/fcmSH
M1mLsR67YicJVCD6nZP76oQUXIeLyoTGz8JAoCLkuA2rloiakldNrh+1QyQAKEnw
d97m/jo8+k5ae1IK3MMF8vOKa8WiVnxXLZScYBpPHKu9CsjfSoeN/nh+LYctbblH
xWhU/2u6m/Ex4YTFGIqQ3rkttKhmxaMrkhYBIUMEW5g98eOnF/KtfeG4kPs/drJl
YfmPTLdSawPpRH+SzQ3NMb0w4mfjGFSnH+ZMkt0Ni2vT/rvAdJIFXtoy5NliYzOw
P9VAu1Lb9Hc6YyR2g9kQHNFPtkeT0QbwaRD7c5o5jvmXXvwDw2NfouqXnX5Frovr
To4zzXsYxfVvQxrsspVxG51QShSw6lQGNS9tokiJvFkBlvgDowI0Gp4T/X/oea7F
0wwhSV1LTDLFDp84b2BHLeYjLGcYWFXK7s6IEmiqBNbfb29XPACs6A+36yNA8ARK
soF+ujRVOu2GNEMDLFptXJ8ruNp0VValHKD1JCvicTZnuMB2vczjUghCOL19C+tv
PH4oAP3G4+e31jDSgiLWoTbSpYOwzRpePfwdQoG+NwIGJtjavIwATz/8lTMpLBa8
kBqAZMDEUJpVUcXoUzG7SB1T/w+U4uGRlBBeKhKJe7QhP/18eZczDiGD69IQeNY9
mII74AEO7ZQdz1cwc7vxslmHzT/1kGp8lBpiYijnX4VH8pn9DDBkEEnineAnM8En
fVke420vgp8UYmQCZvyGOi0OM4Out4At43cH6sk9Eh2zUBSSY9KBdyKTQLbH6JBj
MZheCxfO1R+8V9nTnbdxlGAxzlt+o+fbp0VAbGKcaGS1hVUko/58xVrfeE7sb8AA
63RV7uLNi5DXGBiquIPGP6Na6MsGejAzkQiuCuDzo9Iwe570e+90lXoEXIhpEMhO
ecYdFLoc+XedDFR6+yKWrluS7JYSKn7ygKsGJgkdMb1tZXIqPQOLjNGpIhqOk6FL
KgpZKGS5gKHhMa+YghAUEbfonX657pZCbGBBBqD/1iBvl24B9HC4SbPlwZVnA7sM
Z/ohluUD3ALCrYIbYE7vCuL+oEaQpDX22lYnp3ajwg41jIokYG5M1DFJdItabgiT
EVjBW1bI9+nILBhq3f9q3nH/2MQrXbY68gxcF/2YfNa+HV6iOv8/js63EQYk9HQm
Cm0H1ZM+n+ujMaUX9DEjTlAtqld4Hbf9ThS9Qns2pJbyg1tpt3p3WnTsN8m8U96f
ckS33hs8xAWPfr6vpF+x/ZH03FNNqL7weBMKaYQXkh//B34LyZ5FSSFFu2eXef0k
lmxGcGyd/CnN9NDK18ddLOuGEzuZQltl2m86CzjgIj7y5a8Aj7LBx7n9kGQp6NAr
UnlfyxdtN3ZxSKkgKAeus2PdzjpNkGXr6yy8PMRIq3/Uu3xdXCQt9RUpgPtr1g5J
LtyPKDbV2e2Mf5icOPnTRiL/eX1GDsUkWY2ubLqGiXUuJaBOaxIoFbOU62wc7JIA
vuX/SkzuRe4Zvlc6J3ySb7UcAM2/R6NQMtLiE6mNkNNJDV8zKpX/zOYnhjzBtbKb
cRX6qr13uPKbvAHnFpOf+NrTpc/PgR1bLvgKdNWZFsA3iTRMGqUu8gBWDfuvBIhM
cGlffYqw2q+qAha+S2oCcHcqAS6jaLav0cOLWpkFwJjJS82nGUEFChKJvN4YibtJ
qMMK5TlefyTmStC52yY4N9zc4CckHimDTKjf/pePF3A15ycQYWQMljRAUpHxjr4m
OJIDkGxs6Sxs0yOkJAHymaPskHZeeZZ3Xd+LE27KCu8dEyaQxPRMsce2ZjTqNdPY
un4/xHNQZUhBngN7hrOvuhYGaEcW7WQ+XGBwluicnQtuMIJ+f3MLuUi9pqXfxQWj
gp2zoBSmJfL46m1Qd5r2CaFaxOgeBMv2evawroz7TOIVz+nHTnpyyWxNtroQXcz2
kXhbZx7PlHHHVbZvboqezRBB1msX8VkI7Jp80W98xvw2ZDavBZCLQD2CIbEUxhOH
Nv2w+JO6VYz7uj/nJCv3jHUHeIpDIoW/TVa/s8bAPwerxy5oNPFNrIIXrPgRXC/b
rkd1XneNd1Hrf7GBB0gNOFD3pt1cFqiSQQUNekNlntLZ1405oEqrVVY2mVpf+rF0
Ap3l0VZQt/o8iZ/C5vKlOFvwTfvsPT9tQJIlI39DxG8BTCYvsRD1jSLOOmXJHGve
shfo+yRaaqnuClTcXfSsEFha5WgW6x0njAqgFAO5yIva3asFtPUF7paGPlVxFTO/
jKQ1PYW8jW38O90MWq/cCYBGglVCmFmvLu7O+eoTUv1aMSNauM9H93LRqGqVsljM
eSaF8QTWPCZznISc43WvhJDDtloG6o3tiQjZKwOJ+/XeZ9GAv1XdH7Fl3H77EqqV
fTxbE6C2KFkDep95H21GL/qRMZuCqg9ACXCEUjot5IX1fhk4jT5Oma5waM2Fir9P
G0DhTWWtcH4Uqn7ceu+A44IwTZ6jS4VKJSNd256L5JXweJgT57QChs+CTSnjGwSI
aNq013QixhUQQiPaC6sWg4gzXYSSsT5IQ/K+ei6DMVO1JkHXmvFE1/ICcKfoCkVg
BwQTsWxn0uoL49zcG7Qq5AlCmr1GGdstOXu/+X6AfeTDlUHsMpQZH28rqurUa2nl
qkX1zITXNIcQvJgbkclezNLd9r8elLO87QOtAJ5MfvZEJRxQFunNJc6HCkld1mS+
6Q+ZT4RrW556TOzh6vqASovRovzaM/+pj7/sIj2SFdZ0u5F8livZpAnm5cpfXJP6
oTmSUBmq3wg1m8wTan9gwWPvomb9vzSfKefRnIGiD2of6EHjuI89+zl/wLYLAt9R
q5eOgMGDPrByOAcG4AmwnwvUwfYIfzb2qPUgW3cLt8qDyNEyEFnQI/90zHH9R39a
jJL8scCZC6OL2WTKFavpkTq1SspSABnD/UzCx3+ZR6p9Xf6fgkThKBwsz9xCKkxi
CqtHuv8SivQ391h/vhO1WYlRbC+qzOTtHVK3Ho4OMfP7qDaUuiXGf4quTjSapnik
mbvHYRWX3mjWUS4lIJHuWXJAeaux/WuB5jzb8/dzELCVyaCN5mcgzO6p6nHn1pTh
4AKlyB1Lfk/ue5CHk73WtbzoJnIjxErqsaMyN/5gCilCqNVpKGw8IKX+hevrh1ML
sAkxAw22SX0L9yVtCaebBRiRfZUTgxuPC2ALcD1viVIzKEueaHlnYAgrFcl3tpIL
QMd04ffrRAiJWGp96dlOsTFOdE+EEfHvss8wIILTDuQ4jFsLg9f4E1uk6sHvEn0D
DZpvE5AWZalvRlip6NL40ZT7fvC7yOyNC94MNL3pXueDQl8edd6pgNV4FRIxhNPJ
dpqOWXBRjnf3bmf/+RhK4ScSvfEQ4rgTiqrEnmSHPSRqK3HHf/SArYHD6eDQ6UqI
v4LDzUfvzs5TfdxeZf/0axLKp/vmX6qzGY42Fz1kOAKjnThkjdRgp1pv4EEUpC3l
S2jMiyOY4imnjfPzRJEetrj/YqS7GE0smh8FsFr2XnTK58n3BlCQ74BhVBlY2zEW
WpBmTEqE5Nqt7Aqnch7pGnGU2PI21t+4Oy2F3c7UcuSC6vSLRdxmC9iYLGWWBf5L
BMf4BO4VFL8u0QCy4z3QSUnFbxE82Fv6LfWDxOmroOMaD0dSyeCXmGjcOY93Toa0
bQwkVCoFbu/8+YJpxJWv5fpmMY+fq6egYgJAvESdzT3LW9maxmpPyg9BLbwMq1Jl
agNgVxYkjPwzrZ6SJIb6ftMqM55X8TijOqem0xJsXcbx9mueohIbzBhjFwI9/c2e
511D62AV/Jp/1QKvhv8aqjrSPbDYpOaILnaF8DWuDVI80RY4w/T7BrFe4LDBB2Ge
twjOjje0fyhenI6+Nk56NgDN+Yba4UFv/5yIKKkMt4B/2u7OXIMIPhocxfKJH3f5
gPNSnVbIJ5bq0iP/nqVphLFBGQn7udPP+P4IWlV6yEU8xthXx1vGlk4LFETcFclz
U3z2EerSHepdG/4k+SJGbCPaD2HC2/I/RFJ4MtuWtJ10pZbYXTwF40/CvSvXVP/M
6Mpx0qwtA9QpsdtGOoYw1+hqsa0Z7uh8v3ZyqchJjpsW/vmVi1ZEFwDRl4suDbrn
/EmQC0Gq4NhYlXZsQ0kRjsUnAf38zjIHFpwejnRG4ryMaye4WNEtql299W+cTmX7
y0PXNxB2gPAlRBfu8kbZjUApdndCrmViIfc8PzuaiwwDDnpeFRudVa+sWjLuvyDf
gZpNrTDWGUQZfMTutsXryc54RJ1dVZEAHjTi97LxjICmVPxpU3tCwpDo/MspJJlv
lRtgIFtBbuF2xfyWfJ/irYDbsc3G5XnJNFlr9HyKaqccoYG/esje192cW5/BF+Ks
TkpOLx6XyDbM1BuaSJRlSLKAngv7a+4QgHegTY2Xyf/HCOm3i7rRD3z+0qY5F2/l
1W7sNIUcwsQCEYleg11hxe9UvwMhmIZbOGIUqEGyK6Q+evpGXSq8zRzPgefmGZ8t
y8mjQlcdSmGFqRZzjx5lwiIxoYs/uydcyDlG9zpVSL4BF+4yWkAqMkrFoF5fx1wI
JRK0+OaxCSvZfHobgpy3rzuNaVh/Jr+E4La9Qm7pZqHRVIZiXlLRZINRwR6OhBQ/
zR/H5/p4LbetFr7/xxwImho1SXVFsC16M6S8sq6FNtDOZbUxWiiXpVxKzX1p4Dq4
o6fWYQx9wQ0bEH3l4gq0RjLtN0WWmzTAOERQV8zKZq+9v12YlzuCxk7WKJqmyla1
q8m14W2pHy0wnca9O7Tcn2yExzFW2Zt2a9C366b6U9j4ndWb6x/gpYzeThlaGXk1
U1UC9c8v1V5VuIOOAYNVC7TvXJJCsCgE6WZmSfbe+mX4+wi9rWF2xwxvMExWnroN
OEnEemff45H8W/5mI/RIwgB8jJ/1VlgttbZCsjk/y7XrjQZwOzGJohTLeBHWL+pu
GyyeBm4Rp2exhOX5SbtlNdsvUQwpjnqfDmY+ahxwco3Rv85zqxtd2eTk8LWl5x1W
wqdP+J1xv6zKIBk8DAGXu2k7dZIOdALfKh86gNHM99imCHiS6l2spDEoop/WROg3
pbg1X18XeP6CGC31IF580lw1YfObWxkufNrNtrSjbEbZk4baAZRXsHhVkN6C2QBJ
88jM5YzdGKC3wvYHI8NiTc1VCSqXF+xnJGjXNfs+sVc6f/7KxSGDVyZ7KZv39JTB
03r5f4x6LYtsg3lUrkrKI9BX6KAOBELiLFaewvx0heuyJuQTKJxKdWZoxrDzzV+j
aL/yOjrGWNcEaratIAbm4tBVHq68e6cLMNxxCgabFYHuinoDjPgHrpacUko8R2uB
aLsfiZb+xn48nNh7bv/T0qoxxHkDDwbjsrst2fuPoxCu2xNpgEWcblTgM6K/bm0/
eU6PPYp2IyhM87tUIIOjt9JAwJLJiy2JZ3tMuSAnlufGtKSpzxauv/YdUmJxYGQN
2VR9bVOh37rmysUD3Nm+y5ZfWkZj5Zv0N3tT69gCSr4L53ABhm9dubcE7TxZBfZe
lJEIXFRK2a50PqZcLzeuxL4w2naJcfvN+k94lIGyDn6lF222a5GZsgRdy3W31AbF
6anwjkz77FPabmp2YhOPikZ/04/zNCiU7HX6GbtUOpTDxZ6o5ixwqE+THfgISPor
flW2QeUJuf1qW1xap+67Ep3sclzfwZQJMCori4YHi9C+eTCF+gbBWO/ca7H4diEr
fxeXCmPhpx54xND8HJpeAjeHkrI/4rdYN+RF/Ab/RlAybYztzcWl6qACjwizPKdW
LGgSWycn6YWZiA0h9/u0dbw/XouDV7swvZJz3VtQUXRnhpFQ0ZNzHU0bfp3BfXmN
p03q7chFQ6TxRVAj7log2w5NAWE0lIm+Gu8j355RDNRcIvHDMwti0F7JdaFKrTsE
MX7lxBawM0i6HCTNnuAbnwYapPYNU946RNJFERbCbDaLo1TrW2Y3hyRVAm/koMZj
SVeG+/cL3tJsSavt1kBfyMMfnsBUyA+cmhp5gxwSjFfdMB6xBN6PTKGoDkdDhqKJ
ZyI5nm0AlfJEcMB6K2r4bOicOCKnq7atQlsS6OdyDx1jUcxNHVgMvNFPdkHdj2yn
80cpSjovf6ZAzln3Jdg3WYw0BuRTrKVNU2MMru4kBfA8Q69AnAzOP/lDIBtZOWBV
UdWLMPlxgqO6EB2fl1zcutZ4B0XqgV2+1Ab9ZTj7s1uXrUKjL2px5YU3DTkWKOzV
x3qKXrldjH43n1+E2Nu0seWyJ5AZK+aXDDfHaKWPBSWx3JbDszY33qkuEa7NRfuO
81JvBPcqq/Qpg/UaHkw3BsdqT6lUB2s0ucGFEV6+L9idL9KDzWKp0Mn2nGKeboTP
iZ0a7zPyLHWvALMuCkIPFbkO97fIjxm14gKkzOG+j9V27n7xDtS/F9z7Yzyv/O0D
O/0qIE0T4Tv9CRhM4K1LuME/jEPNvFUM/QLYmTZ1WR7wNjilvP4d+eYW1L1yMDIe
PaPTEBVi4ck7BPSSaB0zxNK0KhI/r57N8UYBXUN6NIdehh4IXuNiqYRMIXnJ2Y7M
4XERw5pEUVUMIyiPa471mVjjHYEIsHbUTxqBdm0ZxvB+HyJ4WSKAlNtdQ4j5MYya
BbW3LWE2sLgqlS+SEi+R2301Q3B9ycY+0N1OU4x7ea6tKBALq1oZsmhdlj4c3hjP
pJADTcaoztQHDyx/u9AUISwhbb0YmXx99ygf6yYqzpPO1FuYRTXuwIvEzGD+VKAg
JKT9QTPxuSW+i8zJrFiFHYaJnGvRj+31C2lhraCmocc+o9Ozfwlixnr+6zT6Mtqe
1lwqqRcB6Ae8BQcbUPWcDLtZ+2GOIYB8kYgMuYMtO3TKZPLBNjMZhgIqxPiOF0/1
6OsU49lzrE7QCCYryvitwmkFxRMFYjcYL4UB0wKsfP6hawICpCB49W3lMIkvtAOJ
vE2VwRI8f3ceGAWu5W0OLzs07dey5IOs8dvq3w+BNZdNVM4aF4MgZJUDnB5RYRVr
vW2eiWdcQx98wX4kWDOdZSypLw5wtvBMRLecOAVfGn73YAuSR5492/LRsTcBL9se
9jExYcGOcHjnlXrDQp6KWo01jxj0a79vGSC2kVp5L6fk6IhRI+F+nZ5CDWZ3tYJk
rvz7sg4ae5pKpFvBwFBCsJU+v8Lh9UkyKYoJvcfKVWd12C44GF6GL8Da45xTVROF
/kIpa4eZ/hBTA7yBBMV4jKUVvlw3A9SyutW5YRE11QG2iltqe5GRk28XoQnAIiq5
qoLemHMnrhce30FVF+7Y7PhCIf/IwnA8U2b4FYuFoflI656fIyu9CTML1uTR44QK
BgTLjPHPo2I+vqw/lSb/oUKWBlg0y5rJUtIbnMIouWTwEazUx24TctevQo6Z7HSj
f/sMqBxL3vOgnx5MGlI2QHQh2tVe0nFCmqrDp8/06kQX6KVH33TjBZbzmwhBx601
d1sd+uZLpKOOIMONqu4ripPoWRcBpi9AFvwg3seqwxUE/Pu9AsctHlNJZdwGA2cg
+0txGguY9Suwup/GobUK+yVYWfhUbCpn9znWpJa6dfZz34DT84ZO3w5dPkd3sf6Y
TSOFUwdk8L27SngTUpJVrJ0t+UEk8bFXNTs5956cES40OiqeqtJHUdrl/4/5SGWb
btti4s2mEdg+3lVDAGjLBDSYj8BOysoVJsJI34DPXFObfC5S2N9CFXYZCG6WRClD
vI6Ar+xmiuyO+ZR4kq6dLDa3M8fdcDGD5Xj4dCkH1Yt64+A99p0Ki5+cpPL6Ofgm
xR8sj/0iXjI/EvdtPzCMcwzz5HkHTfbEt9PtqbbxKbps3C5K8RPIvsblAy0teaXj
ls7yAyFJNFxidMR0wDvdEcEYg0QToWONs18Wtankk52I3wHgHTflP49DRza7b/jB
FsJmPmBwNGPIx5YtrRjwXMNhl9AMdBVpTPDMik9eqYh06c6RNlVRaZQR5znW5qvL
73vo6jhcNnPa+TYSSNebxFlcbsUT06gRkDbnbIK9AJ5UWpINoGzJTF7uTGjCWsvJ
s3Y0kgsK1KUZIz9b0/wl79m7T5GO3czH90xV6zanTVZUHK5LjUhW2k2493qoDzD1
2eZmxCL5gjFpmvCUhRTiiPAOhHdbQxWnDiQN/LVUDYrw9qe1H+G7Etyxxy2rfJbt
SEVLE01NCmy6TQlYS//vST0HCSY/XoO85CdyzN/yXGqn9+i8KEOucoCliGc0sTI2
ioDPdldwDGbSusj+M0ZWjvC5vU0dcHzBD1MDW0UfJKZsC92w4WxZzjB7x/UAtK9I
w8HBPgcrXo+uTRXQ3CgqadYRmXPqWZNlmplQBHmyBTiLiv1ii/McMKjpvZHrmAkf
la6jMFgCYA0A81YJLHrCdQeXsqpbikpBx/h4l6fBu5SS7RCUdNms2YJNRRN3y4FB
KeLN3+PDCXtdAVix098C1Eq2fGnc/AMuKaLnP3GQ34HmmIa6LTaveoRO7uu9e6gN
pt9g5Qj0Gy7JUvJwcVbC7lRKsdMb9nE4Cr2BwX3rUSmZrxBVo+PXyxZungY3RmqP
W2FKR2Pg7HN8fbZbP7jY1NcpedeHnbN8ujbCXl3lZXd9dQBC5/ljEpcUCvn9VFdS
orJo2oqvb06PAnmizYs8LV7CVp/jKzL7GC1SshwaBT6Vtd655wyJBzP21cQtJ2fT
+PpjH4OQ6HITTdZRPex2DETeDcUGPizHc2/LuPrcXmnnLHHYOj7dKFpO5EZAnN2/
P+G8O+SrlZAr4T9469yIW6KwPIOHryll/ESn24GaOvBT5MPgk5O8lrvpQXzUKFn+
eE8KskkzUlDqfoVEU7yLaO7ZZ8MKwEAe/N0jUxxgBPgVadUlhIjTNUvfCHUphTZZ
XRAfMrbRR5dw8JQqOT68snMCVqB2yu5eG5N9sFYV4D9B5rUzUpku71yX/ZgwX+WZ
pH3yFJTeNKOsMqQZbQknfhaQV5QUsXsjA9DryaT+9Uc7NpgVcfXvtqqOM4vnjc31
2bGdb+qI0XKs/KAVtSWgHzQmB083N3TrMbkZM0ZjeF5FLfwCUHwNjqhfRSwHGD5v
BOG60Pr4p+IC6XT8WeJSEDlxkLzkoGGufv2pXePIpWMsYTXS2OPPxYhFlLlx/5cG
9bQpvI/u/mMWlzOiUtCxAXUBwUurfLkCTaFAGFXQ+7U0s6bqAtzuUWB53Jv4ffTy
u8JmUQdPDzPVLFw4nTAUkcBftOWClmpWhRMkOG9U+N79OOw5L9PQRdYfr6XX4HsL
Q5l5Jk99xPKQ0qPeOBRM2x+dmPsgTU9upOWILDcEqzyYvEFmwfxIa7m9QEVp0gAq
uhsdE5GelooV/BS56a1GnDlOBbBLpGYMuYpOb/OTyGCHek8p/cWaBFzZj2vcOOsD
DYnQLYZFN/9vFIwpq5tEfq3Wj3F68Z32+hY82Agtko6nTYLKrDJbg3jdRxupF5vX
/IiCieLtUzdo2s/cskwysuYk5UyuacHx/6WcTUaJIzLhrY8Z3bEV6nx2N/Ey46p5
0DtRxOUG7U0UwmiWR7lCq8jU+PaDHgqvaIfydQCHs7bXdaK1Y7hGOYFtZJUuaI19
qri3itGUmPrwtQSvEuZ0ltxYeiWiPx79HSyWAp5bMO6hUD7PjC6wC6Put1RNZ/E0
xSdatfVYJhNuZmHtGv4ZYJyBHHdtOar5UXItBpurmPa8obcXmwV4ZvrWGloYXY/Q
0IP9IF42nc17eeTZQKDEy22x86dfc+imq39ZKlUJHbEK0jbekAJV9LnWiuRBk7O4
IqoN9ODxploA+owYP0v3l+Po/+F2MQ2ZLLFwiXjo6wSqw7TOuycU255gwgRaYxw3
GuSus2UvMZp/P0mUbbpDUTKhiuGE2H+G66e2MGH+r/jhsM/40/n9lY2JK9nQraMe
XRGHYw638EH5jwNSTNvw/AFBagc3IvUvshe+Twmmuj2RF37TT+zyb04w810z0PLG
Whb3vOIZVvdXEAjjy4FFzDkDHNfBy++RWv30q7auXQjanaTiZhfS/u/XdGDQsUOw
kB5wBm7gee7123IrrkDdEIXOlbZxBSlBaTt4mWrCAO0TWbizmhBFw/OxQ5eOLMCn
jX2CW50RwZzu6QTeZO9fJ+dALLENR5fBwmqlofOBDmKguDHCZnwqS2e70kmiZBG8
0UZL7Re12IX/vzFgEpRYZsdrj0FmkjPwIB2DD7fwzMq5hS83l5ft5yWyEsa5kaLW
JhG6rHmY47KkAGk+U9G+MToE3r+UDZsqQJrkCCnH0NnGizlevNetLGNPut3bkSZC
qKcxCFcCKaC1NQKp2IBIoic6VRWn1VM6gW/M1OpHy/Y+Z5LNX82eSxx2CVVkSKmm
9IedVOjdRCyJst0OddoXo8RyJ5jBO2ZszZqXF7qjIZ1i6ALSpg7ZrvQzCwm4Mk+9
iClvKk9QWrZisNzviJqUAwi+YMeyUFN22by7K2mwQ75xbGdetvFQu3TFnXp1QDqt
DG61U0MZKsx1eC1KGrm3qBtARWUC5ExBOQnQI95chQgUFJ1Rkpm0aPvBlBZpP7Ht
fg/r8W/zf1upPp3XH31fuoD7wiYGw2/3I6Lp0qYpoRZbSmNfWeDtvAq5OKHmB801
JGhdF55JlZjbnfjhE8P3P/QCwwNluiF/+vaigFNYrDQZ3dHNFL0zUWUWl0v7qnnj
G1tHzWpw940Ghu6AqzEZNL6cfe3DvGBqu/VKxA4tF7bLc3W4yiRLvQgBJmuGohTW
L7FUiHElld2/NUNVp5wwB4bpkmNg1FJ7xHsx5JQDZFHGzv+SbuhE7NRpH/JzDXYB
yohaQzvAY/OBN6SX1nUHu+r2DDZsX6dSbnuPe1sI3iUViHWnRFzZAv48mLySO6qv
DZCMChtviHN9fcCB9izPpxiHXTyBGoHTlhKNe0ndSCbB4nyr23z8di3Tw9nMkjEW
2Edk2zQtoasSQPvd+Fsh9LAmytCiJSstKYaBg1wpm3olHasOhi4Au2JQXBHhiBhD
vox0UpS0EC30FnjcqLq0NOT9L1au6nPMCq7pOl5Ao91Tou05Gt1gsljhLelG97RL
MbvUuSlTzWG5sikclq6wrbD80FioHWbIXfgQC3nL40TTo8fhOCzwGWVdCW7XTY45
PhlIAsP9VfxBtODwg1M7tPLYm3vZBITssHli2Dw9QY7dc5PxKc/5W5Dd+FeP6bk9
lDcbtOrwQHOIkLggX2mKHDIAEVD1wUx9L0sUbZFHPpwbOxR7x87TrK6FzE2ekeQd
UQVEoLcu+gj68Sww3OxQlj/q5usQ+3qsdG86BKFZ74e7R4VUmjsNRC8oHQYtyk85
bSka6ffhdzLNR9BC9PBIQfH+DSeG+T0GN3wXZXZyzmNShDwmTSH+8Yydf3gFnJxw
K5qGSqivToGJqhrTuArSjR+2+SPS9QkwJZOTCEPl3oZqmKnYIt0zHe+EOTkAD5TM
sLmKeBxrIldOp3tv49dPSfDh6emC+b9lsbPLsvB+nTvToxJtTNrQLGVdgDcjPuVE
U/St1pDsO3RhEg34N92w6y9qJ9VTmeTgl87/VH+Z9KTEpUj3xBVNVFcpRXZEABXK
FRoTQMSFqJ9jR3AZCK+dTzFIdPXwDtEeVdiAMJK7nlvQ8GFXZ8jPAadJz7oW0aF7
ELVeYcrwy5buwzEXxAPIvkI7rrwzrSWYqoOHEskCRZjdV7bs/jTwgpKU3kz3DY3m
XkVVaqrUzrb2WzRIUFZokuOPd0SraNeP/bZiuy6Tn5ETnGtJB4Ew3ani9kwK9mXG
VmX+yqvNNOcuGTI4IJyvx4pWfNs/kJRtT+UVJ+L6I350yhNEH2WwGcF7Mp7RcIjM
eWL9coNpjTnkLAy99SO8OIsM5XjV5n9RW/jK3d7ijiq56M2SDhRrY8qvi0hoDHwQ
9VCgZodF65dr6DnqlHCXOyHGLgpX9gvap5b7/uki2lSqdaAgv4vNWUt5+7BGT8JL
cOLMR95+XyOxlL+I+hIIj0gJUBHf8mYR/j8h6Q+v5AjaNJ1oYZt2o6tkzRwF+rbm
L5NCtbjqPQ+Lz5PwF1mX0zFwY3cjgA0CTKimz7SfWF4vso7CFUaIJeOgIk177Nla
+9u0R0PHNrWztQMvh3Y8NXLenTPUn7o8PwXso227joXt6T6LvkZlwih7I3wINSpI
Jaq7VGgvdDJHEyNHUZNeI+UMBBa4IYSEEvIzDN7dpctWV/yXEGn/AIcVgJ+rDpoX
2/QSyI77RnJUbNf9hsOquMPGrHjrCwFWWgwCnHw6J5qYZU5TdfkGeMVhKzfSkH+H
G0rRbzOsiXBARDialTUsfTsiyi+RjpiGSMEo72pSQ6hlK7qNCx1L54vmhjKFQ/ty
U/ODZ5T+6VTcWvxSGOfXfHyi9mJQg+fz2+frQ1PLOXsmMXEuok+/PBOVSJRUuLdY
iWuidv7zASatpJq1iMZZ1Hg5PMqG+lFsqm1Vy31nRWH+zzm3F6IAzCAUXZp3DMdx
EQX8xwykyuC9rFrfgi1ZleX98GroJwLzpxE3cESJ8ywFwen/6OMWu2RJxaQ/tUcR
VwyfV8WGus8kF0kQcDiX6Vmu5xudbY9e0DNInZt9x2tHuWU7D2PSnTlah0RW91ON
i6n1GhTwSaIyTeXP6Nf0VpU7M6rhmcXai0bIwUXE7h1IkiVHEUcXhU7S+vP7MP8p
eLfg0L/Qf5eGm3o+jnbF2kMxycltYHl/guHcAtYlrko9n31r2XfMrpk1Ux2Jaby5
7NabhGdf1cuV3Ce0TziVsHcO789gK+UIiOUNrVhT47lXabeSqbhz034/5IN3e4Uv
qtgJcsNHl2rAvu1/nWRcKzdg9w0fkzi0LqJiQ0hQJ+sjCpeEH08AkPs4x6m71guc
ctQGnNoYE+zD0JL6F0y/QIFO9NtcLdl9Srf0oVVOoBT2yfT/WbgNGyzX0Na8nLhR
EXgE/c93k1Froupap7ysKm2HY3T0rGBIaqdtXizYAPY81vem1gnOi/ewntoGlEAR
hZKU6S5uFoQP9wCwRS950EqSNU8txf/rQqSnnXV2ryqyLIZC3or3Gffps0A+eTY+
uIZl4RMMd8mvHgh6DBReN2w9FkHwVKVYaEbzW6A4hNPsHBuVVd4IwEH0EX93tv4T
7gFCmdLF4M5IInVqdvTZjSMo5UpACvHtglR/IQ2jFU0MpL5x77VTPUJ5iKwcOZsS
tV2RwCr9b+ShJQ32aOIIWjx3xbaqiXBvomEO/ZZTiyc2lP/eecNlv/QxIBYJQo9q
aJvhc9GGOrzq1hy9GME7HJMnk4dgEEeI/6f7/dubmYPmHf1QLCP9ZV4S5H/VKBmN
Bqie9uf+19CvYHm0F3pL3VweYNSfNlldK7J75fB2o5z5E/yk1H7xpHjdN0Pp5eTA
n1w216JmHhfXjXkVXjpOcMRo771cZoncnhZHHRp+MF8pz9MgeElhup/kfCKZlamT
o/lr58cVfB5KBIJaaQktYDx2xySTwoJtJ6QJhGrMAFBNztg2HhlLB7jZmDTRQmUW
BJ/i3WDvEAuAe7VIM20MWP3WP1UhY3agh6/GhxMRhC2dXokniFowcejxCGhF8HRY
Axc8B3FuEWW+31OlCSAFYyeE0jgFFtn93ra+7b5FdpASJL/xL5PLyR8FNZ3ML1wb
sblcKLlJffxLVSKRBUZWEdgQgjFnh35ahXOkpW5RvYRCtPywHchZxdmStweiPr8g
SjsfJGnSRBCaW/Cu2iRWV+alEQ7cdgef0ZOMK4q+bWZZsAHCN3x/bVUScBL0TToE
GxV1AO6LUY5OHZWNPTkP+OBUBJdkrpgsAaPwxP8Ox22WjovO8I1OYG0ar7EtpB58
JIt3XU/p6fc5BubX7F4Oy4qVbepj4IoBPro+vRu9x2MG369eGnzTQ8KKx9V1Nzrv
irEAp0SVClbTgG9kxU3/379/eH0WvJEE1zeIiIlnSpmHf8kmN/cWMeQXSremrGuV
5c9+cLq3F1RoCtHtp4PyFueFWRTlK0c961JQpMnUc+va05toG1MslFeBDsIzNRN1
/2YOxIroi6af09GlZtuRYtHQ1S4EsF0sX2vTaAEIbRha3ZI+xFG8G5E2Zv2U8hYW
NdodzCqs1nvRfzkvEQ/6Bml2cOkD9Y18OcDb5R7c1pdNuspX5t3I/AN/ZsPm9sig
IOHeKS6IGlUBk4Ry5xRYq2CSEHSIqkQNuua/Zfhyrv66yL+F2YPgkxgZUr1BU4hb
Q5HEBaG9irAXFPlrS/Sa4RCL0nhvl/bjp6dj4uoR3LRIrMeGxrjlO08AC5LYQ1GJ
mnHyK55Ob4oow6gM75Z6X92hk+ZG3nY4YevnYMbnaHad2P5gHjnbGIyo8D6m1XWH
9TcPFa+FFXDJewpHkSNoZ/aNQ8rNAfolPTnhxub95zMfnRgiqX23+2Ab7CTG5/+J
lqi+Qgk33HQpD2fDUWkymA8gJsNWUhsdI/JiD2TX0Tjj594Un/SSBD5DoyH49Ln4
eqAWbia0vQhmW+TYyIELg7w1f1yYYBORpI/Uy/NrvPRQGkpr8HjFX/Y+ejPBC23F
iDJS2fmiSzHCIs14/Iodv1ajy/L98bUD1avOsFGKHWbfpqidSQNGmdW6tZKjnW+J
UImEFep40bP7Iofl7g2DhxTQrowKir01/BujHO3AUJ0WB2oxTelygtxLMceNSYUT
qupy9GCtLPXwLIJddtAJ5fqeUaXJyTgNKI9YO08ily2vvaTj27o4fc1Gw7u3c7m0
nsyTc6p42p8pGBoY5VfafS6Y+U13STPd2vC29KOjhC1Uirlgf4JzP/XZIX0rj0DV
516sIqFJ/G1gHxF5dn4icSELwvAnQoSbfTdW+lGnLYy68lL4x5tWfwxMtNWGXWiU
Mf7y2ZSV37eoqogrtQQIU7Ri8IKvnLNSPtavf9XhjchLspcCmhqJiTTN6dyCSGxZ
nhXQwwFB0/8LJswXzNWm6cIS2WeS3MchDdQCF3NHijPmyIzKF87Iux4aGxeqIBFR
S+BTVhXyzu8G7bGqxxR2WIWKwcQCZO11aYcyu0tILkoKWUZRLWulEn6BcrCsLySm
AKZuwE+asp7qdeKm9O0UqMr5Gz0jXb6NZBzMT0goo5leBoa92o0qhoakxauU0i1X
EpFFPpqtAw6T68ycDFr3UfI0RuuzUQQFRX9F8qTV3uEtZq99XywvIzPrR7qnTwNl
dlwna7JkpAvLcUfY0S8sJ8l/EYBlFITk1J+mNy2FuXEN3uYmgUJOFeqVmBjGItyR
VT3fxmYNIvQWHyZKKDG9+5gRCVA21LrU5BX3tx4iAQIZ4kw2iDrEzD/evcCE22hd
n80zRsWatV78tCDxtRiuxyNZHipGnOEJdYYXf/qNXcZl6xgv2xIzqrPTl4P41bVn
gje9TAH5P7Xbtvj0CP6jQ/FshFzYTum1NfgaTo/ucmksCKO9F4ZvM1Rc3huVr6CH
DRhD6A5HeBjj/ylcEJrvYM/8w0QkDtnD01rknEE6TZQ9AhGsxlYzRM4J4Fc3DsFP
leHNLVaHNrt72q9Qr3LCVYSeNmFkIkTfxrsn1O3T71JsP17y5MmhRndIL1gn5K83
3anaFFQhtSxcgelsr215aTYSxC5uWlrc0FMK6i95akOVjVX8Z4s5M2tdmyB1IyiF
ak0fT2tgDvAlEjVvpey7bMYOqkvZTf4Y0O3bXJsHntNnB2TFq9/SS8UjgzdLPg52
v4XC3bftWh2o1YKyo83FQ+bJ5fPQ9eGYjUZaA8m3CT8Bj0CUoKeSkAsQ4+hQpJ4V
Z9XAWD394dFppPnynPMNxVhu5XW3rJjPNdYNhc0O/h6VUigNNsliIUHPZ5zk1oBg
QZGqhiNLooRMpkDtvdE5ihVC+bNLQY427yR6xW13HzaqYbmxENoQNOGa/Yhx4bTO
p06YO22cIkDx4HvVq6Z+sXqSuGnH4IJ1qPK+/T5in1ik2NQfP80J51V/7JL+rkDl
1qzrvmcN2BiLbY6kWB/x7GmeLeKuN3sTYouG96e4q1f8c223vjL90UTkAPAtxZJa
pycTTh8+1qFAexO0yIhwdtv/ZxoH4QOKHKMOZ/O80AIH/mVxlwl4qv1SHocJ0f/8
yzAWC4dY6ZTpD3/GWrnEUNCKPo9FughLSg1eb8IbkpQOit0F9+t3Z8x3bnlC8mXF
MaY9EBXJHhj/Iogeyz8/7jyTbrmKzLrl1sTL90vTzpdls8qsbNd5R8R0x4H0m5V7
L6d+Iy+qFaRA+mFQcz5twOSuC2kgmwmozEfmZc+4F2Ld/veizT1AJ7yXSaSpCc1h
gGuSjiHXLj+cvmvfRXZdB6J6IkgMt26xoPy5o8fff1tw9RT7ZAVffs9Sw3EPr2No
QPHWr5u4k4uCT4I5qvLkaGZ/gLajYoL93ye22yGso4zMUIV4+WtFgXxrsCBZc0m9
h+0CEg4M1dhrp7tLQNULZQy+7GlB//JQ8Xq6Mnc17Z0iQ2rjRmAd8p+fo3qZ8ISY
p/sOnti9X+HIn5gDAttTLHkOY2KE3JGxC7soEREwVgXWkkybFdKYRfUjLUobe3uC
D1qZNrj6RarHtgguHe1nQpI05w0ogmWXFAuI1WN1rI3O6I14CoaJQpRKyH4XASwM
tursW2KJScXhffsluKPN/ggvnofMTLcSC/T+IUmZ22zMvRBgPDXjEz1r+mpw+3x1
JciKItA6ExpF0YXBO2nbnuMQobuA5e+jcvOk6olm5R5htw/Pb+dUoWhQSR+8RTtt
tmQfh0mjt93S6W/mUIFu0BHfq99GG7Fv4PMSOiOgH7O6OqaJD/68CIH4ataQAJC9
E6WKUM2g83JOYDM0hDaZJTPyrO0sUypwlBfifTuI96vTZYJUDgbiW8cPdjsmjh8+
K47Y5XZ2XUrcb7hmihgG+drDftQuSgzF9H56KpD6Xw+K8AMCEgAiMzCsCvnmX6TS
nWQ4JB3OD4Mb83wMGfhC8azxBN7w5NejDL5QTW8YeDeeNWmdzCiaVaGX6uYqU7MK
2jQzBnjZG5HI27+xdfCt1h0lK6qvmyi9ZhuiJtLT9Nje4ctz8Pr5HEdyXuJJuX6L
qhgQUu8Qjj7m8W9n86BiDkIg5IdCkLaFWKWa6w2H4F5je6J9B4NBp0sufp4LNAx+
SER4Ejt2QST1Ha+z7jEomoTfags6sVVqB7vf3nVkGn7nBJJjAGUwLc7MLIxA53Ji
cLJnmLWnGQ1ehpoFTBs7GF2RjXK40Jq0ofK34Pue0691NLx2Kb/PJOo9BNTl9A53
31HwJPrtbJFwTiB3pVGzMVHjOxKHTmjrqO6AvsDpZEBz0rhQ8705ZY5wtILtkca+
un9j2KQ58AV2f00Woi8aQapowyfo7F5pB2j8RnhCIVCVaX3tIeGYJ4cY+tj4TdKr
7c/GXr3sTkFrGctHBiLpoVZGY5v+wS7zzTxETfbZ5+0Y8YK5ojAOx7pJVEhjkNom
YV92PSoBEQfQl/aVsOMum7tLMZUwdV+llVL6UaMzFNHgZ7zvkZdAK2p1ZMpl2tQ9
QE2xe50GjrclhIeStvlu7Xpp4JnKJZT94loPj3XfBSxESfULfIQ69GQN9SKr7VCc
vFdmhcs/IY+japEjOlIz7ZEwLNcDFZp1xZgqFUHfueLfmhm40X5y+nhVIhIz8Ogy
cPh7Gr76nyReEdpXN4+0Ytecx2weW+uInAlJcyl3JlqYm3qwW0oDs0KkB8KoXODq
tuupUbMSNgbjFMj9259SoBdve3B7kMD/xMKls4W+0A5m/jlihMeA0o4Fd/f2elIL
vpx9wJaJMEnBKveQgLRAkcvSeJqUkfYm+wCZee6WcA8f69sHe0m95ZkRmgyyWYYn
CYY7gWnWSQj6io7SQnmit46uuxcVFYqYkEWRA69ZE8AekM5ZKISmPPaT0LReX10B
/DU1K7PnqCtwjLwdbWsikixtrcYoLyUtUHS3xGLFgG5WvWa9R7zwVzt+IMgapmnL
OVJgIL9RGbbyBYDAcopO2tBq0+HVc6fTrx9YCOq20HHIIdko8AtbkY23JaxBlIQV
CSZOjPr1ts7hYvgh1OML03hykO3gHgNvIUlZxF47uC1QLJTsrrpUunV3iCA68IWl
z+fpiXFmgwrJC1EkzXXIH6JKD46ylW8DWzQmEH+eE9JkGNZUg472oDy6ZXvQhQx3
Vltn0rV2TCvcbqptsZRJPx9APujYwX4t36oDnSyfWfm/UodiRXzk/oZ3Y55OWj/Y
ZnbLujmRg5iRdVD7MxXAEKXk7cP6CJnx/rjzPg8lBgk4Q9DoNj09KHJW7fiTBRf3
4f3VT//GZFhQ1KdpQ9azDy9wuOH0Ke/rJLDemuED44czKfQuJtm2y44LMlNu3wL1
DdWpXi+78hxsQzHA1mhjxW7anyMVIEktSI4KRkALjtLELbzpw0cH3BRa7Jo7Xp+n
FPXayd7r58zfwDxGkf3RSHo+1PM+G6AxnQRvVdvSFY/tibVp15rSCUG4Ye52cS06
b5ap8abTTvhI9gdjxJ6+pe2cZaEUg3HlfBZErKBuxPzVTe417IgpZ2oeKsKRdMwq
reRA34rXpYWKEsWGssXso8Mxf5N+nH0sDubtpnQ4s9AEpjuSBUikYtxMI6Ifxev2
PbzIs+m6QbbQpBG+G7bOjbM+6VKkOZ+BG4EFRHMFxoeLQHn3JFopkvhBxjcF9XqL
UlOvLqr/WQ8buTQS0ftU6Z9Xmv8yr1gm1sx3cC6y8ZaDwW8L7WUt2aX3kBEY9/5g
VauzswlBTLrlhNJBJFbd6DBeCgXCw/RIU1TbeS+ypxxqkrA7JIZ1RdiBn0OkxcOo
dE2jYbsvyV01bB40HrQczgZQnNz100k5ml5Xt9LSIwaxDF07d8tTsCCGHzCAUc7E
szsZ0ODIKa56t3JynCDcwP3jbpRgHSu6alGpy7dESBV+shMbvZxhbvfNn+6vTSGu
QNDnmPXHxauPBZ8755YsylTUO0eU3yGCfAXg5yoJfscVdhVOlnWLNmBHhLkdDuOv
J1Y8FHsbqB+OCI9vHbPcx2ZaKDInufFavtihiOKhmdkYnXDvPfzuEh7SXOJ7uFPn
d6aIB2Bu93VAJjGVAKVWwU13T5y9KqyYJOTK6jOZnlo0j1suJ9tm27K4awN6vUMF
4kGs7ujWVL7qxn3uGCua6UjSPhyoiknQOMD9todPLW0vtuEoRb9IBR4W8n3IEBeW
0fKZmWUv86ibjjIUp+xAJPBeqppywtDObbX/dipzj4n5cO4555FxEDqSN8kooiWF
AC5Y8Yzp9YnqaCYDABs8qJcnlAtsb+imKDdZwWB3sUNY7eBCEUxQfMDdowUbZJki
vHbrH2LxVZgH4QOEXXXH22Qt464IJyQbtGjdTVw9NViZT0tr+HGcx+tLD38hd0uY
wkroppKFq0o1qZr8f80Zlii5QxQLEtZrySthAIypnvVYFGTzNYugD6cc/DOKq+RE
ZsGO5qE6VW6oulsk53otTWBi/oKvfnehsWrJ8eyquxmliGejNjmAkeZuN8PPi0nR
ii7LZ4tu/oPigzdzKvqKsDaBdPKLtgk80q5b+vERUSoJ2uK7OX23Rv4K0Ai/Mtgd
wg4I0t7aJPIzMyrNNuRK8jsrp8yvYRvp3G3eEgFcYitH53fn6mwcpFxNt/Txi5Sr
r4Uhfa9DidyfY/0w2JRMvk0djxMkzGrLmdWxayVWb5Y99dGVDy14Z9YBUuF4OxLj
04vYJtS4q/eTKG2ITZMaG30wtiDtJcmoX7VTvQjuq6NHRZ8D8I7uycJVfDCgT52a
P21oh9jHPg37mLuQdLo/q1UKvNohp/nCTbxnut/aqrIh1MWcehl02z1VIjkgc809
kcaykNvCq8dfuIByIXE88NOzqCOq+nZKf5rxOfuj6k9rOvY7VVhOufbrmlufPinr
bIDPHx01yP5sP5G7VnHGSoljwS+xT6BUOHdt4v25GsQRhO6Kouc8/j3706itbmYz
z5sf1N+JvxmsvmzU6bipM3gcJEhj98FS/Qg0tXBjy6aeZWLL08O38yQpCV3R21Ze
dG8P/OuCdDRXZZteqmAAOAh6i8VE+tDfLu0eR6XvsDqkvvSBbxaZ4Egd8meBPUc7
3/P+Arv6BSl3SSEPrbzXUF4H+x+QcZKH68q+Di4/o1Fda1dEW91hNgLzqd7LlbwD
xPLQa8YzvdYcx1pzAamujqwWX1JODJYteQRjXRUca0iEiw3sIs8YjatcNVNwidV/
PAQKAUfHY/TwJSO6FqDe5zC3J1X1gr9W8ijwOIUmqAPIcg7e191MGsHoif1DgsY1
u43lE0ZdOGr8JdhFgzXdBhxbLYuqTQkJ50rZe+PPe7lXmtWpRaZtBPst+OC+wcub
y3li5EcOLzVBfNE99dRYOSkUl1OzxPl3tcJt1YpSl+g326Ms/v3FkL819jQTxft6
//PFu0gHrSLs69Q8mPV+9GNtjliNwQp9zm9310xmTvlDzTa47Ribj8v++/AQvM75
NCYRDByzD9h8R7/gVvql6bGJPO1RfakvM16864DbBaEZDehdTI3iye4a6LOpP8pe
AKuZGDIahvt7GeYKiS2ZJOVoHmbxjmpi9egnp8oboh6o3h8SJrHxWAZciT+cv7bb
5BAfcy6KtNdZJMEQlp8gGvp1x/9r0UtCJT4AJt8h8umS8gXJI9dD6woFWNDob0+S
dUDU0YSGfW9NBO0l3CTcGv9P0Ku+PhhpBOyQ6/xDJL0nYyRkRi0L95FnxehRbwEQ
QjAfGPla09HsQLvCSkcLFDMkbCyk0YC7NQC+aMvQQ7FZSqz63BB2mmj1RlB5nH2r
oHrtMja2qpgVk//JQ0PtCQDKETgy6uUSO0UkhOT/dRN7jq0W+nD4yziablhQDI2H
4IVt2LftSvOmmClTJbxOhgrQvzBpMVAwaghiq4itxZAI1GGlEzvlLJClL0aVMS7f
+1rvvVJQGy2eK7RbRIQ37dOwzbor6Op9XVkLw7vYIimUwomL3T018Y+5NR7qrQfT
o2+Dzy13WbjfSnvPJD7U2ZsCsVly4Vu+6KS0wnZ9ZBdqykNk2TrWmtB2bkq3fW7O
niiVPfyCKFrnObkYk1/FwtTHrgXeGXggSeE1B4mjH3PygbdgNEPlKKRaOHT5i1NT
3Fh0ndfbznUwoliKMt5onBK/G90D9bsjGJsaNEFe21CQvzewQek7u+Fctqefqv4h
+T5nzg3LkFv2BrzxssOQyh92qIvwKQ8Xxf0vqGpYIuyQaKiLX2tH9x7I5Pr7yJg9
LS1CQP1Cp9cV65pVlfVoUSCn/bw3dEhb9ncr8TkHipySTL9G2zOnkk+AoBn2x0ko
EKMY67qEZoMd2luySaW2yYLd4WeabQ/NnEshhttEC669kacpvbNvexyPnwT7DDKP
eO8gvYWH47xzJdM1qpm/edvccrKxy1HS9Vu9kIZX2qorUnmEB2xEtol1nuiYXvR7
B1imMycX6c5Zto7866G9Eeb1u/jOK4CE0McRdsjRsYTF9mqktaYf6Cn64LVCIHLK
eT8SuxzavmvQnu1RqKCiTaFXPNiXnobjwmsKWvTwmpsI6HtcJfYMnZ3li4i8qDKB
M0PU2C9zXXO+pgKIwHi0LyJSj0GJhIWwmrVfjGIQ5F3cc2MgEH6tCewaxR88a6By
2vI/I96Zs5wa6MCe7p/SlZHqdfu4WAS4ehPOcfMPhoWhGAfhHL9VN32/c9Yg4Qjo
W0Z+7FJRpqUXIfQqg1FG8/VwKVhH8gEDOqYbjXKdbqCc/+qHQCLAumanQMuARwyk
2sRV2n24jVcpV466ZaU2KAoYAo3e75LGlG81jcnjYAgC4/b1sLo8NNA4dYhESgZU
UZFHPXb0BIAVF9sGIifY0vzg2brSLmcKIxkWaYyV/GkiMOSC7N0TnDz5DZDwhC2l
/t1m1q9ZspO5V9AoKJqrR4ag7K5b5V9Io7t5uzVmBQFUvuSuZfPmW5WUllKT7ZI8
Zd7CL6NnCdp+elSAX/i3fk9NKP8yUMLVdWzG5iv6wSu949UnXNmmm5ptvLpEidBB
gWNmB/GHBMAn5W/33x8M0SWxxxOYPBBLQxotkEwVkoG6+vtjBjBBVFQjvt48OVcI
l5YH6F7CJQzhpgw6qQxGvXTB7WKb3owfAsgM/CQgAtFGqZO8KMHhIKDPEy+ZU3WI
VS8/4hGXWcm4PwKZCit8AJJqCPt8nrbHqeDKaBTSC1+3PCYD9jjsjOgsKDvqFbkW
Rsv2hzGoM55hztikNK2zC+kY7CNVmp8hkQn0AX0BnY6BVsQu4tnkDnwFOVAGN9si
s+qagXz0lbIbQMpPtoDhg8c8SuTfHM3/59uIIotLHoVZAK4YdqQcVWpE2CKknkfA
/ldjaOT85u2sg1WuI6PZpEUGObJ8kCf3x49BjPCXlmAuYMGw2LtoUi2tzBDwJxD/
vUBwaBkWe/5IqhmcxNy3zu/2OAl/2TL3eQwsv0x8bMp2f3J3OGMZj+G+JOMMeq/O
F7/jpOKS3LcVmPprhCadzaamGjQMZCN3CI1D4t/OzyCNMS9IY+SM16kZI6SJQVo+
qTPzPKUoornxN2WW35VkS8kK1+dchzQWRntGu1g6hl28Zjw0UgpNP38qLnhPHmMO
1ZqkpKu+34grPHmCFeAEfa6kgtnd10nTHCqByK7Eejgx7U9R/ChxW7KRmhB66Jvk
3at8WB4On1inAld4f/D/n+A/P9zwTkcHgKZcz3nLmEUh10pdW+NofPvnVQ0J/72v
7IYkcYbsqrfgV4tNP448XFMDup+LX8DLWHMZVbPLfX8qz+UP0WwYoTbuN64hem0g
6+maZS4OKtRqwy3UN+YUXB6cEtgm+Yls9SJlE41cuw24FuKIK2g2vwKq6TUM5tav
JihtB3vDevY5NzCLCWuh0SRBmWU55rKwSlW5HvHAKhExBRet7OWbjYI80jPlEwWg
At8N+55UTUWfj75TyP9NBFuxRfSSfFMicPsl3+Z7kiIwDPKg2b1///iWrP6VoXyH
IUarEmHUySu+/FpihkYnxxW2fUKsjsW14SHLakyD5dvPLRA5vwXVXoV8ETkCkj2V
IT2UHuckyZibA1z1tvKlnxAeHeIImY4xsubNmnoDp6h3R34TS+q+dKM6nnnZknJX
Hq9OQUyus4HIB0FRQthcZEwCVtxPeRp/I++LRKt6s9RYEQRj+K8g/DDpo8eRd9to
PYQ36hMYW9RrS+vGxnsMrD1iwLdX85CE+C2uuJhnvblZQ7LzZ5vKGMECaO2zmx9i
9M2lEpEkHOx0TBXFhDpvLbu2G9nMMUjc1r17fAwRBL7aeUSE3r5G7TM8XMgWs/VG
dsPhA+ZoA+aYrZ1Y++QdQPLPq1hcSkVXa+hEej/6AGgMss3G3NO6WCM6Px0xN9jz
WAy2XWgTQ20i6mS9ENPEzEGWhZxZ0IXx3eKl0Eg0yx2RGbAiYJNYtGHPpP+CPEdV
Yjr5kF6IHnTNWjEghAJGEqbnl/Oi5MssJD9QznygI4rVPQZXKgQaBYXwI9cTgPei
HCZmGP/r1W5n/xOKSHcw0p7iX7aYkxw6i8m8slZXnizzIp3aXirgEF/FNLZlX6u5
EFV9OqtFxrqputcwvX5nf0dNV3f3smPmckXQBuduvA0aJh2y2rgnKlQm6Sl4i4kw
dEUimRgNhaortFsXviXZfqjAqEw4/0UIAHDxZ4uFlEhoe8meBKMhXgpKNqTrpUSr
X4ca9lD7xnll0XKa99qpeYC2cums2MXXO/OxELHCUpNllCbbGRYM/tUba+EWZmVM
abQHaACYWvYrzltlk0ZnEOI6trtJpyux1rLiy9MsXp0Mw7/51/TgD6CRq43bHJFw
WYuNAGPrC9Ra17kH9v46blJTzEtWgK3akO+U/wj/BYoWBp6vLxJXOiA6o/aUz2RR
N2V4vu6vkwhvM9vxihTQeaRtNvy1MuZOCLagjOSlPliFcejUZjgpCaweBaIH/L/4
/Ms61evKGJv+hOoGgm8vCU7iQJtFAQy85MNTTAa+eLd3pJ9QpJYRNOGcq+CYNue3
XZKrFID1x8aFYNikwfJO3JIfoYyMaqPXFMtWI4fCGlK6jeR+11hRbL1b7JQ7P2HL
Muz9HE9ZQwriB+gQorF/LgVebja0uYUQ6CjNJ2nfG454Opb+fB/43sMHkCxgcSUh
weoNRZgIw2R93RydIqV0qu7nZiDSx1cYphuE4tvuWoMdgcZ+X+zdKZJSgro0+n7B
IkCpGfEoA6/628zGN32n+j3rFqdotovt66QctKRlheP5O5nqpc8WVqtLBrji8PxP
3oDmOFAI44QX6rA/dRNP5KuPHSe2TmGbf2bFjqW4BGNTmwPVLdKvltAPHHNlgYs0
3YmP5aWlobkBBROohljHvwaAsBZsDv1xxRNfOQynGb9JQvCsRsuT/ihikXMM5iG1
LP/+RZWqrNy4v9JkSnC2PZW+ykcnSiJJ4UvAmF0O9I1pFzEO4iK6vb7kbad7/FSN
Hez7bxTvvfs0n9dw8zZWyQmkU32BfNpGcKXZodpPZtSVooczXob+CHHn4hFr2bJE
BlLj6dw1YZ5eMixG8eA4NCGctzIashB5xSIbhcEHZwNC2484XujL5sN0LlnlcaDz
cRbEFmAuRUxlH1TJsrkf+9W4q2K6NjAYe4aCWIHgKXF4cn3dwkmU7u6C1Y8tjjHy
BdB5DV3F7T9GpRBiFqGMMYPY7UIRqiosKhLD0h4zasnXxEQkx78+Usg73FOSKQaG
AuPGvhA4CwgtG+wWeLbJcvnOPp6OPFaX8rXQ1vwvsZCZ9EDlvOckzO+8wBCf4rv8
mlsJ8ndljgWr5QkC8ifm1cXNfq6ftS9MKGs5UFZy1v2j2jB0h5fhzDF401UTm8VX
i4UoBBV2M01VyHo4hC6hasP8YA4eFS4OB7AIETUA5Yf+JX30JBbgWZZTnXPdtPY0
o/TTxmroJ+0my2bLD/rcs+w2MwkzaFw3HoKNi0qduYsqaCOcancM54cSuMOxXmy6
gJ1RE3KjpPgCwVQpvBRoVYRypAV67to9SWNdQbi7wD3d20oeXdC4XxN4bnCvBwzK
pQQs6mZqNHRqgmk65YbilF6ZdfPwNR2a8koX/0+tQXSIoAvSffZ0qZOv4QbZTxql
9ddaB3ThbddzoXvVZfb/dXkhxlDEPFxgnwgYulgJS520NUytUlOOu6l4axutZLFg
CjXyn4OS8PSsv5fkJufKnnkIilsw47BXm268OfKqFGNp7nspziHCALw7fhu5JBom
GxrsFnInwbQgn1s0KFe1bTzF7tVeVuHrXSYZLlLEOzEVpShbNiAPY6On2fld9HoI
8rppmucDtcagc6Z2RQFVoEqNO2+ysDl7i5oPIp+6V4jmASg4GHiXUrtPQ2VgV8TR
4bqUfo8UwCzXbKuXUpKnOrTI2FhSyAjXPLBJC/ggZyGnZ5ks0nr70iTjRXKI9waG
kLtHlqPy+JazISkcKVe7+CO5znSxmLzzfKp0gGGkpcTL3qRHVnnjlaCSmI6a8Bvb
A//XMArlgrKcXGYLSHAElEYFbkAfjCcjvb82AQkdX16KX73BbwSNQRo2TBe0DYdm
zHmk+0DBZqCMEtuczi00DqLTusUZh9MEiOv56SpWyLItNr4s5F5Y/ERBrEdjsvzU
JychuSe+QtDJos9bKUQ5fCrboc7qgoehbdl/tPOrnBv0tHYrHn69tiXs7TF+zP6y
w8pNEk52ZYfbP+PSeh0CLFWsflVeXrrkHCH+aUGcWDGYFykfBvdnafinIbIsOepR
RparKb3IQ1jQYjoExnOPJ+ZgsrN8Q7HwoBYmbo/3V9Yxs9ppbuP3qfLaFf1tPlYS
oKjKZVhH6Lei9tWctcdLVwAskQAE+WUaLdDRcIJKPDlBEiOqou0anShJzg3MxpfK
CLeJ2qbRsst/t+vxSsftOOcKOzxServMYpokwrhuwXualh996FYm4friNmkb1diH
8LeqikzaFFcXtK495XI7epZEPWkLxwHVJSC4Sl03a31fXbw1smc3IPAqzlW+kO4G
qN6tITemUQMXjPOdLzIMce0s2cTuwYk8ZELFrf22pkFAFUWUfjR24wKoeiIkCMHX
nuQCnSyXYt1mYVIWeE2KsWooLGe61Blj1Jb3EclCpxiQ+eiLRpDyQYs+34gWkxgy
vUMYCMmwRaQQea/DApEsDpTZnh8bwptHCMigQAB1uBsKW8I4ACHOW6ny3hiwH7Ao
SZB7ypXg4H3BySCcvUj3sIjI86f2rwywMsO9EtKYyfLhOa9/hIUj5uz0HvCC0Kyh
+LuocTePTQ+VUQocbU05twypMeKeadd6rhRnXLgjItqVo6qnnCLGmuhaR8tFHAD0
wcveXIlIJSg2J/C/FCVv/dmVgw9haYXTXpVVb2chimD3rzUkOWm/3Mwdx7eQD/hM
yipUQ6C6UlR38n3Wn5czWFKtQUJqHHbCsCcvXMf3mtphn7K+LhqwdikFaKC07B5d
RZGvWSu4Vc3Vd5eWlX9eoN7eYr+keiw/oJMmP7Uk5g0TfDL+b1BCPIXkyCNehc9q
72gdNoYCOk6HbYFkipJnpozxB1rKNrnHQMK/B5sE2aBvIubnWZ+8CXULdFGbNgsa
QnRtlMAigKIDxr0z38A3JEFIK4MYCFNMcob0YijX617ZJRPfR7O7Q86M3ZJjEXRl
mJvTrVJSSseG6TFsavnZjsF71k7ZFU+V3lJXjKq8wVpdf1AtfPjq853XgWYI2x/A
R1DO+wQyYTHx3eEBfn8L+e/oVjl1PtdLaxK1bZkFeWQewI3/UZb5aPUpqEBYKTAQ
OMUAbKrmnsFmhScd+dt/cKhROUBUCwJr+AjJ13Ayla6KYpyFyv/jAZa+w70eHZ+0
0T477IhQkp+bv67fhJcZyKDQg+bxg1tdQ/xH6jv6efSjRHtj7IsLBQNZ/W7dbLCI
WMsRVw86whYhMaD4demtrde07JbVF3JMWcHEOmyD+OK1dT0tBnsGbR0ullGRnjEJ
QRiRMi8xEXl+7buOtPi19by7PgBPo/Y61skI9KUyCJP/ePVXyaHmxd5KWmooKWfL
VII3IXQ1wPi3cyNxgVH7hfxDs6anU034yG0+MTRkM/JK8wY1ZWm2TYSpjTQKMh8J
ssdKH5+EsAqLiC/9g8CDtF8feGVCKXUUrBBEVs8Ve64Y9d/af5srh/kS2UlHYoz/
q/9tF5Rfi/lkUGwSieq+0Jzhs9XEIb7GeZekVuoQHKFLk4suBoxbzS6ZoKyhSrc0
doIl9XSqjbr8oGqECoNs8oi9wAnQ0kb4kXp4Y3YkFflSfLRkg9nY8S67B5zol21u
L2s8GVuBB2rAjGxOSAAwUDvOAaNExImhP1lg1wNFOIQFYU254WpBOjq8qRlJQ8gr
zpZNJEsbN+zi/Vr2z3LP01KUuWU20oGqY8kLQh2jdDgwvlehICvEdeCLRbna4cx+
oQy3ynmZlmxJT9be2Musu3YYfik145spQlikhGLxdv3j3MVSp7fBbS6DlaxUGH14
vWLiImu9JsU26EYvvzFo+81t/yl4CQ5y+kFUzOEHsKYdOPX0KPUDN404b1YyBNsy
SHxEo/HWRzSSNEjF3onWC6wIA5UZu30fDa3+OXkL4afYH3l8s8dzOAL343ViitM+
AjyE9Wau3FOaoppOZ/hjjTwwERctS3xbA2twx+HGxaVm2vXuOhTHpu49J3tOXkqT
cOnA2IycySTStOgRPwqm+IZhgaRbHpnASjZeW4yPUVn5wg1Z7sNQLaMosaaYj7vw
ai+EebRbhRWUcZrO02pbOh/Az0YSvodywXMsVMhW8eAUkUdtlAhLTyyd1ZdSfjFb
kvym3YuliMdVeRr8Y8/CAjILLNgvJMlF1EakGmXi4FHLwqc87hw3HsJhNLxsTSLK
bRZY7Km1XJd9Yuug3ZKfcASUwvXo00h9KRkaVLl6Xhyn/qXFnPswMg8WIr0GG0iA
xFI4GqGvFdRqrbSNBixe/QXfVfOIRXEDE7xjYLMjTNhYJwGDlwMe+hgW/Og+rD5F
Dc6biY3xC6cPYpTY8Jcvm7OLz103RC+3IScDTKyQpFT0JZkqOvSl2yfiOKHgomTf
8svcOGRYAOeFYad0slgIzXZbSAc2VJYOSlwmcG6WmLDz22sjYKH2DHjZErDIau8e
Ps9IFqjyYnwPPM1+Q4cReesJaCiXzcWfFw5rgQVPwoaZV/xc27a828F1x5lyMBIt
jzEN9RqcZBwm1cpP9Y2LIfoYxkjphzNBhMBSZ1x8W/cOry1qOgO5H5Qcec0jCKfi
IUfGv2CYW5We1DcSRDu14Acawx8k9QFv+6zgKpDQfg87PebC5VQnuHm9XRCPindx
qIp9KwEK6V8bDadUHC7NBSR1lGtnQ38hjtV3c/l0BLOwJ4W5GcFP6pAny8r5Yq3r
s5Oj1W4a+H6U3W2SEfTwvtgdVtX7k/uvZMC2HLbePiqTQV8fpufeNiZFyxexRQSJ
rd6ci3wy3YnW8CvpKPr9Jt/OkKIikzpBxMjOqW3Vgp8XbgvuUeTZg1bOzGag0/m1
QcDSGAdBvzUaGXrEVXUna9ynPbfjUAtPdK8ikPOD/rNay6mlzwcPXZ96sm5mTFv/
By0413EOu/xY4fVdLozZRpcdUgzyKyitW6DK+peKJp/+r0ROaYX/dgkyCe4yOwIz
BkLblgs5s6wXh3y4EjhqmbqY10IFrvVdLZ4u5ftQUy46W03rUuAXKHNi1JQ7dTfB
h1He/3sJP4UhUDMtGt7y93SDmXNvcDLQcWGgXHsuFlSICoRf5panbIVgsOa4RLrH
hB/NwKuau2+NUCutSPbNKeXJT1O3F2KrCx3EDC2Vs1RU1knjWOfoNWjW9mcaJ3B+
azU3HdJfH+0YqibDM7dvip6ehTLqmsido2stB3fovC5Q+OQsIoMpxfCtCW0NuZ62
Qxv7nUuVgc7L1srg5efxhZHbPJ8ICC/v1Jf2Rf55pxVZbiDNJEEh6TqOpu640Zdr
kYl42Fw/6yFdzYf2xM3LlO/Zzq4ZhW1saMxcPH9J+O/DVoXu8Od6bKX2EeB4R70x
3O54pHIsOp+mRFhjtHw5GyynwUlgbh5PA7BGwzqt8Al/FzjclX0RYYK55/drA7cy
/wBfXsY8yp4TYbME239goeGFAvnoLojTucOqASDicX8+DkDjbA7lGcYkm2fk31Gg
WkNpmTU+F0mYn6TLK58f05YP93gs/Blq0wfIVs2lITtkGkrsu+4VuzqKpfI3Yovc
hXRCjyyILI0OPZBEkJ/lbPboT5wdsXAdwysZ/D9jjjOvdT7UOYn9clnBba82qk5a
BC7D/zBHzY+1mb9QtcAB9JfF1jQSn9QY0/f+LAzl6AnTSzj7S5VzRM+teGODbWHV
2OAFJIp4+i0wwpb6lD6+CXQWVbPEKFts/BgrwoaWoSIYmeu+AkjW0fmVBMKCJWtE
8LQFXhMvwGemxj+ocNrh4YGLnn31YCnkQlUa3gLNIJNjf3r7lc0yWuSpMlWL6zaC
/LNGeF7Ysjf7vkY4Tlv9BjgoifUeCqmumnu38awp8X5lO6Wu/+/MINGCJCjhmig2
FYRaYSuiMZf6HzG5Y8j98mOI2QUHk2LK+7D1w9gmvSo=
//pragma protect end_data_block
//pragma protect digest_block
6XJrLK1n2B+cOcxBQJWmqa3ybeM=
//pragma protect end_digest_block
//pragma protect end_protected
