//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
AcUmxIXbDGZdpLrnaMopalJPn0btb4rk73eOOC8+A9bPnghnbuukMa5ysylgcyJz
8X7OLVErdYOW9mLcwKFsn9XBorQBrsRbaM7WhCUt6knCoJzmgPFmqtLaxVqy8Vlz
/mPGjxZtVLb2KLdF1gbEag9ru16QWRiORI3ViViGzc8twKZQ+F6Iig==
//pragma protect end_key_block
//pragma protect digest_block
70vdGhlyAl+P/5ulAMsy+O3oiWk=
//pragma protect end_digest_block
//pragma protect data_block
HUTQYaLOAjQt6ELgTvam6NVF108dZKcraLi7P27Jv7Uva0OZ0CDTmPxat6gyK0Mt
sXk7akODc11FkthG8VZq3VBifNo/zTniBXZ59kG9C8dgMt5ZSDYp9uTd+/tFRdnm
7JXq72NUJWG3FLFhEKgFy8tqFjA6vRuDwQAVv2+GAa2ddzt5JM5T4bzGAEFBZPf/
kh4anJfSECVgimxFoc/3VBHhtXIpIBb4ae4xg4KEI2BDDh1yZDONqe9oRPtp3YdD
R8G3Cvl1cEzWw1Mn909fqh6pT9f5QwRYN+/P5urFgrWqPxA/9Wf7w3ur3tmR3u1u
nfGZzQTcLxcM/ucmQNntjdTbaC8wfo3PVS4jWLOOpOgj3fyuPoysvuMp1kbqmC6I
oLsIS/spkw+84YzIxldEDCrd+njo25+L2yAqq9NfbypTRxgBbeJhv5tjV3eBOHXl
ci/2BeoB0SDBz9fUUc7g8L2mSeCE3TMgaYv2TE51Z9bJnNW0+ZSrtmg+hEf6zMuP
OlWpEXWGRu0m+9vk9tV2736A6d5y2xsnqCMAp0VlinrHYhjoI+s6RjjlkixsPh5Q
mIq4OlMUWxHFKc/PRkuSlCzzK9DGFMvEBt0kDAmsiYrK3L6YZD0JLzU89PZkp4gG
sEpCEacrUb7BMhKsHO7CNbWLY0Z5+dRXYtL/DrXk2NQUCErC9lUfoDYAkYar3Y2F
Cu6IezBKlxQXHTQpKgGw9uzJOVhBjfFvh+WYSPg6kUYhrhdi2JkTTTuU7fAYFMUA
VqWrluODMDiVFsRDRfjNhtWSQqs7YLMhzA7XN3kA303HSD3HZd/JoKPQ4h+MNc8I
oGfQW3FuvHjoewNDjoE4OtJeNof5K7T7hSXLlVW9+SXYWf5uspINLuX/KBqYUSQ3
LQwpo04M041owBnbA9z+ubXPGNoLA7HtguggoR3iHJ/kL5BMJBn5lYrBzLSuLyt0
BccD+d16yN867HxkYt+qA2sMO6LgWOuQDoekHV8T9efUKe2ChWy75TZWPZR3UL1o
RJIAKqbbJBhdOWLR6JiNklfzgYsGbmVaJtKQpwTzQ3+YHeyrF3SHAx24138jLoqy
gV46hl+DwnoQlAf+i3qd9OVtffNR6Dvg6FjHhpq6SfLIlydDcJWuWKZzCXn897UV
Xcm3MhjKtPGFj2Jg/xliLk/W/CgfKyC1hRYS1n7o5jbxy3sejzhX6Ktw9pnL7NfW
h8Ux0ym4oHIZfBH9z4TmgP34Tra4NNmEW7YFH8dpV+3n4LwCA/QFtLwSQdw4Sdfj
Xi96oCjfFpWAm/wQ6ukIlwkSFW7TM/pwDBfoI5b+Zj/pKWMK5wNDYLu09oPRdtmj
7hj0Eyo7HsBBcoa1aq464D0Vthg4GuFhjF7iG/MvGEMT25tS83Il86kZnJZWYCuB
TXVQE+t6o8/wj/QvZu4cRcgoYw1OaYAuwTPJs491kxni1BAt3ghiGQb+Ood8UOa5
JvknLtGL+wyN1/h59sJq5u6VzT0SNcSNS1HdRI0e2lX/Lh4gPv++abUL9z9Ve0VV
Q/bgfd8MSNlB9wiv+UU00UEN/Jdgua3uZE37wrnx5KAbZeisYj1SxpE0lZ3p9ZD/
3tB74+ONEd65R9krEQ2qTCTkcvkCXmTEoMm5qJET1OvsErwuYQ3T9b/tYjScRqKf
x6xNJxjYrqoi0Yi4982OG31AvuiGLZwpcJt52HuUz1Lr+v9jqkHmvEc96jAF/nwJ
IR+RlwVgcB6dSr4qmQu9QwO4ALUOr8E4fGCBydTnSZgo03nH4g+dxTKkA/V1KDb8
ukRUfSvPKoceOCxwRx1XSXHjEk1PZ9gb+o5GQtGymz1A/rxKse2fQ5/YzmC0CvRt
Nb/avFZr9NcSVmAlHtaQrnowgESrrmDQLy9ZGHNv62xCShxmLwG1HH/tVcNjEkDc
SL4mSrETeU7Eanzrzxi7S4cxfBfKUEItFsMZUyizJ0sK+JGY50I+M6hyHxTlhJct
60mAaglErrtWeMb9+hWRmyVZEylNeWCcQUXgqITrAU4d+GFpyMw9TRA6zthjqnKF
sSzSkw1x4JaPBM/M5cicEehBCbbMmQ47TNtMLXjWBhQ/vQqigE9b7eZ9b7KdDt86
DXB3eTfPRQhpgSrFNPdB9YItFVhjqJ0qP7Kt9jpZPTI0axxJhtepso3p9+1aus2O
Gb865I1oU8e5ZWm/Kdw2SHoUVUCBlHs1Q4+lGoYj5PhsBkopT3DMeMRKObI+mJRL
xZBFzpKokJYoueuyK98hmNV7SGJ+4TTfmFqpgFlSDb5k0vo6LsuPWVlxjylUtxx3
JLZJ1s/aQAiBW4edkREKAXZeAee7eWCJH0lVJD5HlPcpaWlJ8J/4QGbLhBld5dFE
1KD4ioDf2wbnlZv9mcYs0VWQ8gtBaEknRv1XyoCbI3elpUIeSOJHzG2dxBzC7Anh
QiXsJfk7/73JDGg3MuWj/vlgKAs6TDpLeIWeWOP6r3m11C1FMAalVf8Zf1vzLV83
8tk360Kd3MLmACZZ2VOKqvUPtIlGkS6RRd0es8D5+ftxPaL0dwBIUGaIKic4d0W+
W/27s5IVxJQKlyljTdsn4aWAJGSt1Y9QjnsQAl7/0sNJLQieYfu76UE2xiwYLRhu
k7w3vqzyrkk9+Ny2WodeVg3U2N7Uu9CWtNgluK4m5V1/5SGFMxjSmHjxiZvfCccT
/uW48AAEJfagZD/A9M9CxB+njfZGkdA7EQVqX3wJ+gFLpSpprOUZ2lTKsRt1T3m8
vEe2yea7ll2ZwctQT3x1wwI4ISbvpYL6L9w/skDWN68cncAl0iu/t6uERvqn4E7U
bF6tsoB70a8fgsADmJXJvD6xdiI9dgPck1lUQuRMzoiUxNGewsQxMvdhT5Zhn2QG
9gE6KxmHmceBoA3K9iQoaY6doLDbdX5LzpNmzw2sk8+DxEpXhpOgnfb8v8rDIo4z
Hoz+BEc47rfNj9hHpoD2/EQGfSCHSQj9QqauUwidBqnX1zbSSFMmod9gMplzCjLC
iE6tUBr8B0hYSen9OjjW3cDPqaBPIT5Ubc+sPrRS5vYeooZ2f0dtDk5lr9RsbyEf
b0YdbW56tea57r/2/FFAGUFm5SO+0X32i42h5+lHSbBJ4KrRJahy4BAKP2i1nHyR
nf4xu+bdMiTDLMXuM8qETHXzgOeyUzwksVIjjAhr5JMO3YdLTBLSw4JU3jpAc+Y8
b3AE8yi5kD/2V691+BhlaTQzIJDFhNBqAxIwVMlEFbUKCJ0mHt60+xZpvNzq8dW9
wR2EjiBHhfzw7C6fzc5gLiAcwpxPZOVNTUunYcmoIdK3mQDaozL1mmVeldCbtjYl
sY8kx8P3tiLwx6S8S/GbyOrq0YY93i+c2dsJ8UrQJD43KvDHx4GjOdRtjiJAXz1P
fnVpnY85T+PKx62aSD9mlHg7yFx80bjJVxhQyUmHWh9ZR6WmDGTveLOQSkbnqV2a
yN32bmb9oh9VqMvBNBC7XAhwG/zL5VJ3uSOBU70lpRF8mE6nPg1FzXmPIidArIoq
+OdedBtJyfFK8r7qcfLq58Wp91st6wL2gmOrEpuZIuLfUWsu7orhe2KmYoxJOzhR
jaA9gbh+lsuL3sl46W3LfRk/Y9q/BYkTrB72vxcIiake8qxcYcqDa4uMFDc1UCWr
2qJ2hSJoAqLLH+qmlrg79UNp2TvInEh3UvpNQWlCTUJJLVoRQ6X7vx1c5GCeGgMA
YthY0wUMIduimty4VhVeDgX0K0kFb3fYz1zxLmQr/w8J2aCDhPyhHjyX4dBOueYT
cEY8Lp2blntv2ZC8XDS9pDRKf93PEOc+rpV6YDtt9nR+NkSixRpUJh5P9N9jjYnD
JvUFb3131jRfRn+YU4WWW9/bhcXd2mVFGycZ4L7oa8SQT/8Ea/KYSJ18YdbQrTlp
98fH69AIrmRTcCqldbMcKZpSurGhU5WPvQsWpFtRI065ka69SLzwCaFaDYvtMnrm
V+2yNTH8AoilZsIQX9DVrCimDaAjfbbd3drjnSzKz3piX8vS8y4bF4odajjJEeTD
UcwnPN8xIrJvWEpSxocOHf/xhixRhIC2pDvV5pG7PbkC5u8qk25w5ePd13v647FT
CUtTY7SaHEjbnLr6eXA5DwA9Mfr9Ul+46RhtOp/KCc7XGmlf/amlCJluD1QAtqAw
nCXZPoJwDd2/AQPxBGuAKhw7z58dazhqVe7lhhs7IoJdTeClvuYA1HBrZFbMutOG
46vz53mPijujnmPyDCihKhWuAhnvWIegdNJdaaSl4TppdYco1Yuh8QkkQvH2nCky
mC7zqMGqG72qdcrmKdEwlYEN9eSzhFbwMBvRVhr5Re82oEK1CeFa76oxQdtG+tRt
KC+Z4djU3mLQedSv7goLOoKkHQQ0vzuYBM4HDSlnjQKDncJD8BQeqYs5ELqODc5w
w3eqTULmo51jQK6AaNETn+NI30VYB742eQPESGX7weH9qcQhsH2u1vFjZRcUDTEt
7MJ/vo2+aKejTrsQznSDKSREl/ui397X3EvJSKCT6PHwuOYuSatPUmi7ovZrhGLL
nvgR5RidwMudgMxAetzhwiCYap527qGhy7nJadt3UkPu9ht2EiMPbG51MofuXOrF
kjLa9MrJjbh0SJECxC0JzHcUdSVGMfRdYSSGIMqyT65mpbTwt+fDQfOnUkq9GINB
L4M0dmkgXMcx+lqCk1cDKmFBzCADFdEIooLZ+HbIO0f6prX68FG4Gkmsz/fAr/XQ
8mNAAqUXdYOiK7p1vuXOkdxdb70Svm3yhNnGQ5GRgxYvBeW2sxK5v149cIxHVVuA
/b3D6y4gau3LzunFTBmiqpGcqQ2NmNCHXKv8VfGvQt4E1at316p7tUd/AqWm35rV
LoH/HgGgixt42j354orOZitHwse14MZ1DSuMjpNYj/RMZfGKZiEjwEg80DMb2BbH
rKBjEhLPKdW8slEZIDgt7556Z2q+34N3NLxMShFGEiFt6TC0b9Xp24Mwt6HpbeBF
YAhiz71FEfbAZqsShdzaQ4RK0PJQ7hp2t2aLeaNrtPrA+VsKDSc0eV79uQWG813K
v2nw8oi0PFiP/Xs30cBucxhFPShgOAJ0CX8qpDWrXM0e02LGPF09png718SWXv9v
2t0uF1TkMviPozIuBmqvZaakwJjmhjTxKqJ9pDs2swT4CaDpW/YhpoRTZLkrkrUi
+x8GhozzrjrCdFRzFsBkxhG5iNsrFqK0uEeM1A8sjteu9SbMwzL9JBL01K8xwG/3
hS7yO3jkSH/D+UvQBRvAz3k+KfQFZ+0AeSbqI4b99JK7dymDB1Y1LFkcgWDTqmKj
cd9VoaU9dVH9RJDDR+Az5dOBA0orHD3NJfXUcAP0bVO8m3qscFVo08jOUZOwO6/f
SoRHbF3Qs9mC4rOSloZpaEtyXtDiZLsI4t7ezGqm23LVjMtQRX3bdCTQPue20QPj
s7kqWkCY36lP51Qis161jEcMv5cfeXiuvcinf+jtaZuFuKU5ICu0q2Xjby9iFbuN
/+k7BKOG9mTUQYgH3Vm2n7JG+zkjZ0AGvJq6Gy4ZVPMxnkApVLNm/3r0KVjC8QJb
QSkuf0GA/nt+L4NqXM1DPiwJsxeas81xR7qPVfZ2yJ/c2N3h3erk4W7up6Afj2QF
0rVV/8oH1ds/uSziRmCzhU5hzTggep4QVhoSl4PMjGzyuvcsU8r/9nCklf0N24s4
rvWB0Ppumh9aAW6qCjIr1uQ59rLUv6xcBZyN/Vm4yRJkQWYFy495lruAXtHr1ZYT
dZBs7NJpHt+7ynxtsAG9e0Ac4jcO3u4Vq9+eMExC+/goP6csP2hNWbd9tGd6MwFQ
+vfTfrvMewR19GzdmRoPyb8RjnapXEfX3QvOt1EQxNRjjR7hj6oEv6N9V+VrAhP1
7zh6FwY7e9z8X0AGjpcmvS/0pyOmRaVLz+ROsHaZvTLOTAW28YAhZp2iTbhAGQ2V
FEgn5iDYAPIqmGgFcbsuzj5CUdyqkE7+Xwrd5vznwpBEyUytZRV3RhJk1s2WcovI
g5VA43CF3pIx27dDr+72/22te64sOr8ZwZCGMPlrbS5bN+CjorJliD4VsZDKCew3
yc2O2wMCZohi6sqHZ6RyCyLM9KGV7M+Ua2j/kFYsKYS2geO1y7j3IzW4zrL1WKtP
2PZAA2mxG2na/stJkpbEVSk8V/XQ6as6/2MLLGgHLQEoDpdGGdQs9ffDMM+nq49s
gvMbkAqnEVgoGs9h37vz0fKp90JYikZqyQOBZGZ6+fczXC7zG7rZ0q9uI+MriFj7
qNQZGYJ5kzZpprdy4ANjqxP6VmXkDf7OlxyQHbxAcYx/a5xvAC9vvb5iIxN5oPEr
zkIyH+p5WyecEEKLfYvT3cRpKkJU7K62ri1BFBOeheG1x5RoRvsXI6jurZ/as75d
z3rf9oOvUHzrGEQ1F+JQ9tHbIiGh9qPFexKw6LrCUH/RLr3p0JHAd6O68IONbrar
CL12dYN2rbhufVrgWdHC2AcFiqx0KJLgAZcbSP0tNaQ83zaekWBxEnKk25uV0ROS
duqDulbAJU4oOPPxQmT77Efdyv+xA42l6vYahuveia1xhINeN5LgzXEZ+tyBvlQ9
WAvzkkQz4IoE5yVGoRrS1lHw69SXyoQ8gYoLYxgN5Qw0LPAdHER7LY8Cze0EOXz8
lEkF4ZdwZGDtYQbAcBOEtlnLyr/1EH/SZd/MkUUneDzz9zUJqqEXNGmHl2dwD+nY
NfVsnFFdQbKlTmDZLRaypm61Als9BkJmVFQkHRBWWrb4DVqyJGh8dxwBUAfu+5jZ
lXypotNHqWeYabq1kX2jJ8mKx14MMYQDKEZx8+STcDydZTkw2hXisLP1x/8hh3CI
IHtc7PmOKO/HgihQ6rel98Sj1MbNIPzFUZJulK2WQSpmHx4EDmoQ61eWWOEwqPS1
nUCs5VeuIzMDpVsb3iiy3a4E3aLaB/UIgmtmQb1vn1dS9wUySnkhn+ATusThUpU1
r2lmLdEMzhSBVDJTClRqUDLGQBLEuL5Iy/xhWJXb0wDXVMmRpAvSMWOiPGqUq7Kj
sIRImN+4NxGeJ52A20cEc4P34f7IacAYxqyQVPqF5BShaPyUYOBpmo+3F68eP2qn
0UUphGu249ccJmH+clhBBblb9FdpCJBBe/XsI+E9XP1BxYszNrSqcDBboVhp+O1l
05y4XH12pH+nFmtTUxVTUbX3zcIpRq1K4nQzQ+eP5MKEd8wIrjsuZmA46fb3UTnO
ZvLM/LYU6Jqey4reomzYH1F2jKGTvzIWdH5qltAiNVYq/qyN+sSr5t4Hsvfzrvkd
Kls6t5cStYI7vD9Ggy7pN7xkFTp+QOuJGSqdP4neeIOZXonJnUwUyV8KY2zNOpi7
vbfWw8/gaSQjUT7hvMSmLLNCjt7TZVPKwryaxYz8fJ3GoADy0uVozuls3QAJklkP
JGCNNdG6Lko95VfplngJqh2qaoha2+ZcFdoY11pJKJIcRaDmH5DEQibkp8PuIR22
gwk8q1UzJImdJqPsCjPVNM6frdpeQyZw35g11t0lurVg4XStxeXRmdhyefoESlsT
IZVz6GoVd20MbjIvlKo/3drgjxWbkikwklrmjSyIZyXWP/RmYwIGh+YqbwJeFqlC
/b3PJOf0N6CiNk3wfJRZhlvEV1xrdLWiUFLcIrhhnqY9D4/w3DQ2On+WLrHf9k2/
FjDojkD1avdx4IDdsIY0JsuxgMnQ1y+fWCMclIllEQq93RJwfMvPXOOnqSsRox6M
7J6D6pAk6waT7cx7MbHpIy1LAY5DoRwz83/A3HcqasAqsPcqaw+Hi5MxCScf7TWY
TB3rqclM7bb9u9T/0T7H1thm+FvdzFQVHXRhSZyzCPvwRmxszZZIYlJwchiaeHiD
6G/eOiut6uEZPyqAeCTZBz5xTspevR2IN054q8iM4AT8fP+oYd7XkN9r6mkWkRMG
gSkY8mLLvYrPk23iTtMI4ppD+AGxBm9DhK5gcuNCEb5EO+Ka1MOF7IbbpDJJCuCJ
3+CB6nqMrjRyqz56po5iHWkjIwooNUyebuMXFFLNLqxmxKoQ54kRjVYOPFhNJ5fW
xpQArPtMA8nZMbWfKBZg/b4WFJn5tUOFGX8OSkvrmR8qtg2RzVVFW95byEL4Dxem
B4rtWZFDk0Efr0tSMxOUyPMlKjfebLijH4GHniRFyhq6CZW1pzbJrZ2JwodXOAnF
9KgpMjaXauBkuz8v7mbybtxbpA63BMxYken5jEIS7I3sOoAfVJRQCXtk8iFud+MM
zl7yNN/gTw036QEm0/5HGU0KXPkTqIG8lxq0w6M+E5GLKKUBrNYj+NUcnxcDs6xg
2XWZUBz1AesWetXXG5OAlcIbLY6ytNnu9A0VZVlOWFiQytQ8DjeaIenEl6wiF4ST
QjHNvy4vgt2LM0nooOZz4Rij+YB8YBUu4pRANXi3gleSb8e5p50thppZVfS5aB0M
YfOq79ARTVYHc2Qc3YiJC/d2qL1bWHaNVizZXMZhrJKGGdv6pA7i54WeK1ppqvXT
Hm0dqeNH8TsgZmqMWMsio+OmmQ1cXfdQhbwuBjQwd4edsbsSRXin6AFvqwsv5afH
Rkh4Ux4exnA/Sj6QM1/+TDdGvXdQuRwObkoYbLbP451d4/S8nL793U7R4ZCwP57A
nMboSckVUGzLQJDCuwOEq2tXj2XU7jN84BqduVI6/fgrs3UzszqpP9zqo1bVOogD
zdSbiScxsO9HqrZ94osjTsMyTNvyho2veGvSkkbwScaY4HAXd7oPd+wqeWCa5sXD
6PQ6SoW3/tdd3PqccJExmXXmRdD3ZyJ72ynggYK71m57QZyDmP7ka76YfS1RW2dW
t1v6tdFdWBjvxLAAP+46ziZnh3H4LP3rmibLFeHNNC/fgbL379C4MwMT6XCVKCR2
keJOAvn8q4ksagXjfEyhBMD6GZiQAoCvj/jzP96nK2SJVzhGl8q9Z13JhFFY1KtU
BIEOIDisCnIAXdQFj3wY+6iEGWFi2DmAIL9T5TH7KAIikmJzgdjjDBY9Z5E41VdO
gflhewr8eSwdnf4M95OV0iq7CreittTaDwC+uv9PSA4WA+Jkjh8NN8zgoIW8kahE
qRh4ondGZFqEA3ZnSpZRV5EdQLXmOFGpOdImkUxhlTZ5u5X12znoI5FVd1N99wxZ
ozNTxv44ZBj+OKuMffopPWS6PE0sCSXTUG5ysiXosvsULDD65f5gzmrWfUAKxC5l
XKTzP/IJH3AV1bzLDG6ZQ37RxKbDqOkUGnH3R2dM4ehkV/akrrwpreUewHMlVwzy
8S9WpFifpuVc05hvwQzH89LhG+eqTzGZxt01hOUTmLN4oCQSfseiqYNfhHqHN35c
VYZ6LIHiiSTpXRdZh904BgyDEgaBQIloledKE4Au4t08DuldA1tZrDuZHvD+RZ0H
b/GurUUpms1G+7Qya8IXOFJt/vhwhjWBgvJotr1zngNuABQjE6Qob9BiGVS/quvH
o14RKKXVNcMdjN/9YL3cY5mhavCq/7fw/3+5/l91ddcTEDs+LIZEoU/pSG07FQFx
vVJjyjdCXuYjOqUM5a8MbrNOpO4ypplkZPV48KNOXXkc7tI04knw9SvwJ1dH0/IT
6AVZJdtcLej5xVyshtX1oOa+fP57TkeJYDPNTqP9KzwU1Iiz8/k+rCoSBX77Gubt
by4XVWOalvbZj16HyLObRKd6SSpScS4R+NwI/WFNog1DbZhtBraybk8mcRlqHbNI
72K0DrN6aN4O6egFvZYa/+piiUzNRTCqN9hkz3uRfKIst86hH875qJ9veUMKsP/b
BTWXn82tqeKrBIqszA0lW62ICXeo2iR9RRP7W8mlg75k1hLXa1+jvq2WsS6YzOb0
a4jqu9UW6mo1cYWZEQo4sHwOdTDB15KOv4zP6pvC67S+0nW3RWmBeXEnEh2b7VdY
jIfxz5pNJ6Oy/HxKUW71BOQQ3eGJD++HFhrl9pHe7RhIFWgnb08E/QrIiNkaF8LW
Ae0Wk+PiQo0Ur/FJLG9X7zmzGUbn2e6kXJ6bkNiO/WRpNe1bwlciRqeE78Pf33l2
rI3AJBtTW6nNFMzj1xP8+w1MUH3gzToDSiX8FUFtigx4dyTYZuN5SSDRXINFhOGx
E0gV4zMWGece46ia8yzsovmAMFSYtcfYp4wynG9Kjbl5Mm1MZLlaLePR71RzQ9Wc
XPtBORjRTHabMCkPH1XhPN2YWUvNeEvs2MSvX9OhlYrZfk5fSf2NpbFuDa6ai1zf
jHyX15io+qrDx8agQv/e/lLwu49fxbzRVavysIFvfR8M37xqwfBp4j9+vqrh6sTR
T6GZpeFKGjns6wLzW+87noE2pYmSGkf9tfOGBoddX5FzFkMn3VkfMuXYpvgiM2ND
nqC/SBmr2Q5tGyk3pFlzlzGIayRRWLLo6GNYTDygmDSWw0B0Rv3XiCVujbHwrWAZ
UWPfOHp3wHBX3eRl/Musop/JsAKp0ODlN3cByAqOBL14/lmh6UeMRsGgI3rjZVIQ
34qIfAyjs5hh33Z5i/rDxwDjf8q4/RSat5zZoMMsOM4hNFTpdnqvGumJfDn8WFHg
wWVQ67DLGfct/oMsYMcq1UEr24MwMTYldB2kfyAtXZBomw1HpI0uJ65aZdGPgBzT
8JgKlAGkSKsrNHvwIUJB7jHA7IKwVujSfNy7NxXqoResbhox28DiBizTHH1QBR0z
CGB0c1xc7pwcjUxEzQVh5pJOXW6v/1tMKZc+EGZhY6hLDZ3NCj20fJ0kSEGmeWEG
1dYLBwet/pieweH2d1RfT6ScpZrwj0g7vvM5KbMiAdHs+/iJ5M2mwCe7W0WPTtSm
jKRuk07806a+IlovMz7sjbKQMrmvPjdJBmQEIKSSTHp5bdugi9hiooSqfpNn7gnF
xTBQ/6EepIrW4cvUpXMWwXgLmqqPSN9rpgdG6B5p54eDugv2Xfak24d2PZy81Ytn
icxYB/dRwDFJ4wNswa53JfuBSASDMf39s2SXi9f6eiHEQGKwPhKLR05aZTAvRfuP
PRmO0rNfGMbgDAwDp8vCimjONeJ+Yt5MrwQwTRFP/AkmwOnqyN1vbw2UcGfowTEH
ZM6/ZEdELiCwlDvXX3/sflVIVHJ/ssIdAZEmO0pn25Ifd8ututLoC8X5NWALn9Vy
zkFYeFbg1Hh6OzgfjyU4HeEl804snHCtdJGZVZEj33LmolNcaP/zJiK4IR3ozTWD
8gAwTG986+pLE4viMP9nrSp+KuCIEGERw3VXER/XYGZ7CjKZL9J467IU/lbL270z
srn1Lj/JHGRhatGXcgTrUyK2zaaAubxr5R0Bu4Cj4T8PurBgIxHjdN3pYTebokUJ
oebFMN2d9QEdH5cYuSpiHTp5cD9i4VF+JjzRMHLPgXBGTc75FjdJ9McM+z6UtCKQ
z+lhVnWMW04fbSUqjouWL+qbzzTKfhduvBXoFRCKbTEg3DkpntKTRyhic6e+gHzE
EQJ/PvBLOeB3SL8rnniKHeSFAm4z94upcMGyCFLOICbzwpA44l2JPV6ki/0Jbs0c
pc+TcghCvQ3mYH06Vkw5/cKGdfcc5qj8HZWLGJwACzZbtxaNIsPEvILZpF8dC/Ks
kCtzbRmk/P6FdTHbyqinKcbTuS000c4s9zA/E/Nsj79jdWbZrE0rddeTsdOqPn2Z
Ktz7mdmZsB4BI9fEBlYci+2UfBoZZ7k98tlOjcq63sezyC6hOi3MdtgN54qTZAYb
BukiVqyukAIsgGHbs0ODpoLaUPl44HWlD74ObZXU0mpTFYJeOnXS8/zBoUCaskrI
LHb+o6ZDw3P4z1JPqW2dytCDaEsMez0KE9ECXb35DTbLKUZCeSMZ7eP5j2vXzSzw
RxgEeKLTMnvof59x/dbxYXf+dJQA0ThpEWVy4appoRrDwGr0r2cbSjHYcSmhlcMO
4YDN97dieM0/9vvLT/IPWF3DKcz/zXWkJtyvNwiMOr6lAuVuVU0hyNGQAfKfwcQR
KlJjauWYXoo6g151utU4tBMcoVhCsRfPw5kW2q51vebb9Yp/dieb1sMh4dZ0+pcn
sfNjUbiSoaLO+YGtrrdOk0/JGFe2KYKj6LAxruyFyUZ0bC5t+uYaKFk6ihIUL6pC
fHF3UdnaX9KCneGRFRLtUsre2LreGbRIdRCRk8AkmHByHaL+vS6HKg3zIQz1n3RQ
bonHx6v/QhqLdu8019j6Y7D5Oru1uAO6Q1/0lkhsXw36SF1fq87LSPP6yHTzzOcX
MuM/GiCAlJTRFcyR9ugiKsyQ2L1zryJ6MeEYM8eGY4WX3+H2PzlqejiUrczSmd+F
66OLK8vxCo15Ge7n8J1xMdAej3totlXc/1S3B9py+/6yk79I3LAjKIyOPYToyQDx
POVFWaLHBu4/HetldxARXWczeQZbvdZqvqEgYyt22ys/aoDitIXSXV6KcshUEgzv
hj0SJwUvaUSr3nOHJ+gNMbL3nCkSmA5GT4g9+PN88RMFjtZuS3+WRmCPEYa0ERjQ
WasHEe+YRBopVs6HD+rHpsijtewZEwonME2zm/IXW+8wWxHeh+D1vTjXxtR4tt3V
9B3x6pXNXnKrbkAHnQ0oZL1f4Jo6leHAOQaK8EZahLwdkYAdKR0q82eLuVwIZEmx
8Yrpj0hxRrGrOpNe1S1covjhCIN2G26hW6NvTLWKiyCesvQwNQMBcdw1/vZpAzIm
kGrCcb3SUCNNXMDd/hSoHeMmMjq+ZPOGRZ6kyYPz6q7yEx32Fp2k7FUJ+plMCZW7
bQKr5s5FJSAjWxRKYVUxJyMYItZMitSeG3JmcUeHHwH19keluH7KpFbP04MnX7Bz
dwFWVl9Q/8QXQDehMrD3I+Igi+9eb4znhFrtDpW/iGxz8c8dG/EILkAbH2JHfg2e
akwtzVtsJmvu+7+v4oq88R7O1jENJ2LWTrC60V0PuKhQ4AwhOJpOeK3B6jYfk1O4
ILbwriSnUpBhCK2KPmbxuFx0VRgnILS5DcdmRNWqY2alhnaTvfQWItB82Ooabp2/
JvW5P6v/U4hIYPZxj54JOEjC2fVkq81Xj5twElW2KlEnckSlPOF4bpnrLgZWduEE
aLt+ZTQmYxLx7LpoAI+YzVSaxrpVqPrzkD1rotsDI8n2DHyV/foxMsy4zo2sKo1Z
MlEqqCbo/4jaKVCePXXb65IedFwO1Erc72r9jMb9NaFB3qSQ02LylJfIHZc0hIms
1RQ8HxROmixBwo/PvBcEevbl80H/r+o7Q4N61xpxl6NoLsABsqjivHKsQijCzvJA
xjYRHw/grhoTBQ39bSzC5wziJlSlrX3Jctoz94AKHMi0IgfAYE4enmfPs2DP2XbV
+I4WdgYaS91CqEzO7jtUxHYvYjx7zXjFGYt3Au8NT9wheCAzQf5Op3F+oE67O2Ra
F/XbCI7fD+khyE8iaXE9xqryk4Mu79ZBW35+m3BE1Kv3vgMBEQRj8/Z8A0wOy1z5
wmoC5DVMAtPS0iUHA1DakjUbFMGmr1kF/xOzNWUvwvRkXC12six+OPyS2Fm2OrHX
KgiTAGw8Ss3n6UmjVSTE+BAVuMa8DgNovc9Vqxr1XOe8k9SNRaDWh7/TKnhnjego
6bRoyo+4EqKr/U/Y+y8isB8WAKKj3WeB6E1ghaQ6HhtNcygvtykuVaouDiMVKI+s
zBSHmsVHBkFQ+s5CJFALY/YsZAlFTm5+0RESF4XsCXbPLuAJ17gYUU5jjFfIDcBH
YVR6MP2vqYArPKNpoHik72YnHc/dWe9Jf7o8LWWuh/s6O+L8tFAcyQeZMcyC284h
2+p8KrxKqBP6eqnlAtuJURI3T4jJa0kTN0ZqFm2d47CifeI5zIkY0GmTQyZ3dG/U
Lrlalz4TUOUQ5MJ3B2KCnzINY/5eVHOHf2e66YYINT47TEGw5BUA8GrroDMXeWC+
kks4v6+fDJxPA/hAX5n8XzxKrc8RvVhawogG/NnRa7TnSIXmLrI5m1+zI6gskgfd
3/5oTzrKftZLxA+9CTO3H9+kn+5B0s1zBXTE54Q9wYuMARQHoxxpVjomb4NVGX3i
frGkGVw8Bz1tBzdCyOg8+dWlybEvoYiUcfzj3we1mh1HpkmGFH+cCBWblQINiSoy
jIIsWkjV0Rv37pVkxLxtrvqdevxmCnS/NSjj0zXTnaciUqqw9eAw8GK440tmuyG7
qyYo+/rO3pa+4bXtqa3+q5wg6NhvT4t8LjPbguNCYaCKadjJFTMXqPRasDCAIcPx
f+/JBzKIoPwbI/bt79t86HmDHl3qF92pUiReFlH+hk9MHylI7ATPt6Wvr6jxIkJ2
ULdM7xJvQl9EYMU85NcRGgruMPmtsRXNtjzyChgHFht8E3htwPntuw52LI56d00l
isDbgq8xF/e4xlxHvLrGb5UmTAlyG39N4zdRBALNDqAZE6eylN9BEZqttopYcyLy
hGIH58QfY8sGK7IW68aCvJY6PZqt2wkvpboTTnNFUq6fkTx4D7dCFjh1gx3ReRqg
llO/KPntvu7ChlK/HBrT8yEamiIGPeqq+Jtd7mZHJ+4lVUZ52oeulHLTb29/70CX
kIaIl0bBtpo5URKMKg0whm715eXH2fQW+2fjAiGqBm1Xove7CwEeHXhnFPonQBv2
iTliXXxARai2bKhMUvIr38xFZP554b4da6TpAwnJTS0jVojm8zbzQKOk75lmZphU
WZvVP6xUMeZAOTeK75W8ZYWwd2Kes+cB5XbtOhMqzTGCoUHvKLMI8/7l5yz7isDJ
aRbJjIWAe3QPuoL5iJZEOMb3ucdspYbXwRUoxhMEndcbxJ93f9RbL7ZZv/u2Kxww
GgowD1HX21AJLLLm6YlztN1B5LOSdTKmV9hTXCQjMHGQqGPQaVh78+5x8huYz4e1
FPA7G0bnMkukvugBLoByPcdjb08HJhnsZfGOsRJvN0E7NWiwNpgoxegxROYvoypn
OxUG7aOguaACesZoiRRTzJgLYoX6czhZgGvK0sMb7tphTBWVvdU94mvjBKdSnuvo
W4O3AfrckCZ2LuYEquB4EAMPQ9HKpFU2YIYyaIChxK7dxwUCUrKmWK0znmQuFL9t
ZyLVgZl4gquj4EnFS01MH31neKZLmhfsZEqDNlK45DgYXrwLBcTa1Ttbn6QSu41C
n7AEGa2sEEM+lBG+RcJM8vNfuUcGwIVCE/olnOPnTmcgrIrRXH5AgyM08Md5bZ1t
01t6ECU84toWvmvBU2WPNiSTYEQNapqZgfVUEIBUE2eqwEHdjDxT2CGzufj08vGu
1jM5sJ4lh7RYij6/FsDKF7a34Z90eIYSsvExexrPNcI8Xd7W3NUStfqs7HwZ/0oA
S73TU9CMocqOwJ9zUlVZOGmBIt/lLGiiKREDuz6MpVzZcMoN6kCqFYIRknMnJQNW
uK3AECvoCiUUwbpIE/+J/gCmk8759faO9Qefev0H8GhL52uDSuXpWa+wkg9IbR4r
lJA2UdqGOsz1sKoDv1qRLFl/KrsKVnCvm2+u/zNKina1+LYDvyfjw9U6o66aWgpa
0aq2OeXJjcAN9BSjaU7JTJy868LQbi9nFrz9mOLmJq+b/7aRFTOLEm0mgmbEfghG
L0k9IKC0SqtRiBS8Ofxhnb0HzEIEF+zmlrimECVcZccUS5ORdj/tdXUT0mxVcVTy
H/sE6N1Ce6leZqb6B1embssMhGYFhXXO1hsOMIJW9eTKU8mt/HuRzhKIaXr+lhAa
oKdsVjDJI/atMvivXH9UhgMiL5lt4kp9sIrNN7JTCXW4JWK37/mj64Cz/rdCOVdQ
C1vzwcJp0AlxC/oLaPos6p1ZvP6sEfNhMq3Fl7zNSp1o0edadLzaShXlxE8FHkWG
WUXzCBH2czAYfoFiw9/DwnQMkjEEJEPgbER+8OKHIX81+3Z5fpKIOYVrscCn8b2H
Et6mXhKfkaeKZBHzZ9N/U+hmuYxleiXTPI6VrPJT9BXwynZQnu/jLmBxr+S5sqcW
2vNilnjS0vLvAHVn0pngzjRFHcxwAvsZE5/ZOUKYPSROvC+FhpM1C5cgUYPctT5w
4tCV5JoTs5jkp/WnhfW8rtGIecXtpFhIkKaG9jgr+rVPzICUKJRSeIue6bUtVkJR
YeehKZI31MoQ7mAQljTBdhb08HjtygOvyyDDPiTDrvDnrzdi+DeyyoDUt9P6EIIC
VdAxA9GPWFIL1pjFkiaq3UapOaKEpOot9nXcGGxDx3L0p16Nhxg/WtTz6qGjTNyA
rwIByZMJrOs6eVe646XssQHo6XR9KWboIf+c5N+OXoEYisHWW8++UgN1yU3K7kUI
d3jllELbvKwBa25MbELwoMOSAvXVxLvWQij7PoKYIhTlU174+5F+jBLqyzv5vcle
q69rO5hmb/Cbbol8zzDNwSZyu8CvLNXcww3sFm5v2fqzaouwthOFH3Nmpu8j0nN/
0naUnBfbkfk33rp3D7UhhkCXzNtgQEMz1848rntDFs2bgG5HxoUaVpM69vuu6ap1
wA/0zAI4gyRfiymHsOm7G5qD3+YFRjDHNxQja3DGhMxkJwDK2vwMty75qUfSDVNB
NfGNj7fTewMwOEvW3u4fExvnYk9Rox6hTjvSTSbuskRgOrwfb1gqlWSla+cE2EV4
M7XhIXdyZd2lEV9uzNrbXUCEb7ZZpf7qXEmSqeldq1+eRMRV1qxEmxyd6vPECUTz
0or8rIkNhNBu+OTT4ou+2TuE44tUXNhea0yQ1p2iRCYHZlTcROn/xQpf4jwF5NeG
oKj7MR49iIuUuRJWKjGwmnl01yJBA+yajuVqsNYuKi8daX0vsi7GO3pYdGHcfoj/
5JvdxkgvRtO3OO2KdnnXQorjEYTaBtUYDbabURMeX0gBp0rlbYe23A1z94GHO0JB
MPA+bhTXazPRrNs/6MHGdisZpyJbq3iZi4nJxvvI+CAjMvzcabT+BMyQ3UqBcjtr
DaY05PUAO8c8KADNDNnFE3ohgoe9YzQWMiaYUdkg+IhZIrrb+ISDpNNyx6pDkHwL
xSO3vi8jRvvIuGzaZ0/4DbgECzsNzSZuV8iSGLt9KEhK7ECa488dhuOOO6yvCmLh
zIM3JlO2gbh4fHWulLzyZqYnZ4+ELhikZpFViCsai9u9iJMIElvCVGyR1h3+zj8Y
KBIKSHFcQ5TAMQ7WspERzeO0HG0S3VctNaOIhh8Mnucbytfowe2kpBB2QmH/7ZV6
5ZkEmjBqXjLTDb/p6n4HMitkQPkwKZDILaG9x+KH0oHEMuPhO2q4gk5EIf4L1gzJ
GDOT0you+XpZAhAVyah3umBON8oRL2JImzwUlLkzcwwrBHBrWxDCVRaSl8JjUo9d
g9mvexu5JVU5pg/M740RJHW5OGc8Uq1FdZAGGwmbZDVpqn27ZDUHG1akCUuvqZGW
FKMO6/4J6gnDGU6v9c3Xsv9LSuqaVCJaVEYI4aR73HaxPR1u/QTM3Mr8R3BFDhD/
OJdlHhbHulBTRllevpnSs+ez194KjWAfnKtMV4EFsUu7kJsdVo4Y1KBrHoIyEwDc
fVVztUZIpxUr1CnE3S0pj0I+en8CL3iSK23A0ee/9Ag+WEqivd1lPntC+9bDnbkt
bm6c6pffewmKM+sy4NhsvYwSv3NG2Wk57PsN/zFaVOkOxm3/Qaw+sNIhfDmu8/d1
2FZrSDuAvIL/wpQC+0UByXQd37EWak2r5gcbuEE1nQYnItWk23mAj+TJDGAG+V/R
wn2eCKKYyKKeQfm+yLsnRSO1hmWLyC/aLERlhDEKean8AyQ9N7v6Z7VgdvWeBZd5
FWaShLiVVXidg0miBPZHb7aoA8DHN0bbfSlCzoa5cNrhJJaMZoPtON2Z4Ll4w/QI
FtDnCC2Be6ewfExEb7ElmWNphl8twH5TvKWACVXB1NqOd+3rOFSggjKV3FnISyMJ
j0HNkRI3LemXlUS21BThFSOMHkgs9EsqI1bKnGFK4YnIvO2/8Z+lAaCVVUKtQNhE
pnpKZdlhu7bR9IIvb4RO2PrRSMOJ/0eoncjN/KsTtVWXsAYh15LrqvG2dOTb6HPq
BDHiq3SOEVMUDems3FmNmMzliNWmvAScHqNy5XAEfezRtD9ffoEto0pRqSo9beKs
qRIuY1kE0rPD1NyPpLiPLKzKCWvMi5wlQWmRgdOgTo7G43c3yb3OqX+k/8hVRF7i
hr/aV2KCpKpk4Cdl0RQIg4dD5m/0+Off8bqbkwY32556S3EIf7ZOZYS6C76RE/Eg
5HDxE9A2x8lxfi5U9BOWzuFNShkrDWz5rkvLrrVO2fuRYcTQ/y62H7DCt9VSmIc4
9Mkz8Mdy6VGioAwQM2PMKwXpYoGjsV4GU5aAP/+jh8JSNF3wjOoITEU+pRXSOzL6
4n0IW2XjlPpb/ijRMvNdurgwztepVhLu9PLe8VCx0YlI6wsii0O4YCDIvSYphypD
xN7F3i4mDuDayBQ/S3JS3Otb8SEM4zBEpSNDbbtgBq+Eu8ATbskq1efutbTu7pgV
kwXI8wlD/XF12m/qIQqkCmk0A+6/u91ZTFXv9bhqOY2S5tIqOTkuti78CAn80MOG
uHCRUqyEC1L1O2bT8t5hV81o3YTRUw/xkODf2JeeGjahln8hbfot4bZYAL7/N3u5
83Tv7+0k/6e/oH7PN1BmqGXJkFz4Vj1vXSAInSB3DMQXpZUVxDu46bvNVJRv7eV3
i2HNp4SS63/eaeUEmf21eqK98kbf5YwisiIvoEWE700JnpPU/9rsfLCG4vAppEpk
eu3sLns82e5nxhLIwJsq6+ob50VbMyDnS+MWLM+PcQGB3QmVfVS4UBTZBSCoaXos
5rQqe2UJXV+m7+k5fdZJgtan66m4gIUrxUDn7yCiX6NP5LFRPu3cjxZupk0IfQ0z
EDUWMtUS2rkfyhzM4IiQTnKYnVyOnRsWQ8bR2cN/F6UuXBAhYJbJfPLkjQcr3GpT
33oaP8M/F2FzQyotBz3hVb6cSOW3LOIaJupO+dW4GRfNqrIBj01btb+gboB+VpVb
IwbzFvHOUe8aL8Yq6KJXCvcSXkAhW3fa1g8RnxwSkUy1YIr5DPYSFasIsUc9tCxm
0zVKSpNscA5wEmNZHzIOjNQI2IIA/b0BuXe1r2/X2Ht3sKB0+JCPKnFgR8lc8n4E
8NiveExqYx3it6hI7c88NNf5XOX7PBT6xDPfVcJcNQQtRQTbn4NTijm9Bt2OS0e5
kR78wk2JyBEq6ulRvHokorg95q/BD6q5gDmjX7emV3izHexZtkiLD3dg0C1+SGf+
f2JIcGQuI/9o+S/6nLXDlU54b+j6ALHWHH0abudHps7dYLAbes27HfEq3GytjaJv
RKZ1FutI+fJNlREZKVzHWG8a/WfDvk2SehNL1/hhIqqg4JxQQBVzSMkkyH26pLNv
el6wONWOhrZUEGfUOarB5uRjlfoYyX4gE26qAOFai2MTAW6FfA5t6pupnQVSkpvK
XDc1kpn5Adt4R0TNf1YuB8EHbWRrbWXBr4ZJx6935kEzUKiC6aw/hXEhL/bJ3fzU
fgXr26Cc1rJYwWEDxbS04+G+qmXNsSq5c+qb5R4BqKtbJQMz9trjBqYEgjQxOf5J
dIpS4Bk0GZytSn014RHJl/G9Y44+cwGiTbo3iw/dfJTr37jZ0vgyFAsYDy4TFyvh
p+hn9zFpXTjzILqwRX0M2IOuA/cFFwcK2PeITDxOdJYxUKriqcevHkqlAMq2saRV
ip+EL3pvbr7oUdy8zSrm+lMsYK5aL97lrog/Tuc2BH+25aSAzDs/vWXd1zxM6bkb
/7zmYnF7vlKgrcREyuXvWURNBuc7E1s8JgjaXSYzuzGL8bTUmuxNtUXuMDuynGcC
YpXzAwjg2iQsZQtEURd7qET008sbJ15uvVgo8B6CtXHIzi8pkjJsmUzKAZjHwvts
2h9GNRD5E26GR7Zww/lE7sswt0xD4Qz0n7plgiN9NQryG8dtBUcmV/yGsLIgsSn5
PK4BeicuDU0LXEw9lUNDJ66+7KEAGfTYlIT28k7gyMVPqxnofpWkGOTU4svULmX1
sUzZtsotxFOx1uDTXYHbIM7TWcBru5ghIMrv/4UDTcibRwZgHq5A8Fq52UAJk1LT
C63PKU0BRwtgtsj88KM4ddF51b8V/fLVzxTY9CIRADksqPDZJ1fg/fiaSbZ6HS1L
5HXXZVvL5o+VTbrsADpbWPRssb1HNhhARGyvpSmjQNg6GXffpUSoGKKkUz9XZKUG
bEMP0mCexer9KGNaQ0YagzfLo4vVbLHdIIRWHOtPnFUAKo7c1fDfseIOWDXLdyeM
Bhrg2voRnOHxwydgYvNUJRTG1Ev7Qx9ljffR5LW6e5iyWANqoi7y3oATtSRk1zfI
ZJpV7ma9YV1prDp/xUq00mtEGHs4R5/rnYXzRgQcidVQRjEHWaVxr/rGxSMbWvf9
DmExhTkfxBS+b8/D/3N4PZNytOXFfZgwCiX4aw7p+PcOKwGcZiP1aCT9eVFPE4tR
bUbNGFyOW1K7riWRRXV9lQYCwcmmuoiNnKMBlL6xl1Cwbb9HdX9cyeaSTvVGsG+Q
RHFtdFw1xzJzowtpGTbIAaMoh8fnw0zBP8co/wijBeWX0RcDTUOYO/CsmhsOTxGk
L6NKknt9sXxg8uy6iH9vC0ctk098B5L03iRxQIUNCoraTx+GYdM7K1aA0nMepH9y
K1vvYNHJJJV2PkvUb5RgqWuCDEYJGJ1XhcnfS0IT2Ngk0TSGoNcOCEEbaB7Eo5Bu
GxTKZSxI+vZCbIuB6GcqFW4ON2RzrmzJllayEkNPUFvzpUNzHNjGwwxbwf7Dw0z4
wSNExm/fmQsw7nawM2wR3MdZGBmxilBE7XFRfbLS+aZH2HmiMUKokRJZ41haYmEH
Aq8pPo2nN5JuQGYOTvRJeP2mfu98wemyRm4lv3zE+AdGqOfZW52taQ4WV6dmxoeQ
1yVAvi+1OjUvu17BB5pjuoCjNW+19Hx5euQk6uAyfK9WMDDcHZDjbmEfuzdFU/54
0MGYbnH+IO3Q0ALu6PbQDhe66wqfNZLwCNXFs8aX3dfw7PJdOPSJXBEZyPya1FO8
FLY4m3IPgAEIwIiCi/nK2oRwJB0zZOyA5ICOqUZ94D/ZkPv2mu3/25Q1eXHlc+np
pZJM/bv8FJ7Volre4IFY5jHyCwsye8tSOKbv2LT+rIgLxBJSMLZVOQANimHT/yzn
oN9SzJCC58z/XAQ86AbHdPm+wSz2K7UYoSVVpW506XHxnhqwIeS8dY0Q9Q1XwaJ3
tA1xegC8lwrDMFBRvZaOIT27x/CC9wr53hv8kc+QRaFBvZm3UuOGc2Qlc9q5rOls
jwh/zif8sW5ieDmHlSPB3UkiYn6wz1tVarxAwWeMrKKMh14fNeVkuU7/ENX2NUtc
uB/Wl1C4wEn00WbRoitHxfANsLfk4hUGIh7G/W/jzsFZRcF9+1ZOkXtGoMMdSLXs
uodTjtYzrn9wrxFIeSvVde3GrBXclgjHRiE+akzQ5O2y0Zmpul3xJxclcyqFCPLn
VKtjDq/VpoEy0M2mUhjiRZ6CfT/sgxM8abaqVdLpRgPbmAryZtERN4wQMTqk2sMJ
nEQP8QCVvuO8mp2VBzSPj/GJULqxHvwxXyABlM0IQlu7QQZ6ZFNgmtnIUFmJluk2
An4QsJs6BJK97Hq1uN/cz5co5TVDfPow4bFGRc0bbmmGC7xJlwZrLu0wHt1Ww0bE
1UtNl/itUIq9EB2IJuuu5EXQ8dztANguueUKwnQnrTKl8BqJEIRF9wZ+Dry6WJhi
N+Jp0mbkc/LaYzw07RzHnzoyrn645hc6SbMlt02rh8ta2iqcLH0CN6j5239XsoZ0
YaBhxlssU7jUR0U84HNvdxYUrMC3pwcXNoKdS+ALqMNRUuSuR8Cuwh7Sho2C6veX
rsK03IdRj9WxirODFpTxNwuikI5L9hwxMeBnwy9N3eEquoUPwu3EGUQrpzVqreTP
q7F0W8ftRxRmi4E2chOkOjDN5ROUBZSDvGDeV1vY6ZtVivkEYKWgg6Gbsv2vcmPl
Eg/v37jcxuaFskIR+ml5REp0oRbZczNCqcbtCRB/jl5Gm+Ju5IsIV+MWAGGsHp5C
NZvO6hX+e7sbNi78FF5aUrHfQysaoPMFV3JOTetqX2jCki8I2gSjf9qdgxeLJI0M
vvl4JGq+VJEVBq0XmtExbvfvYaX9sMWdhvJxwopZxvFGp7TC87zOX9UnnvqNqwnJ
Nj/v4UnkRcU5eO4mPxYjlgg/ME8XMg7PZO11VkK7rVKKMgsSBmIJRx+QRp3/udXK
+1HSluHBUMeoHNrpxCteVPI1m1UnPQYEo1L+wzPai4g5PXDxKcQvbIibRA/xY5gq
rhPE7C0Qoen0ExCcNR30MY9RzCXDQsx+6uVOmazREYPQqTLhlu+YmdUqiyJIUzgB
89wk5DP5YQaElY5C6ax9U2z9wf2ZUaoq3dW4I8kHiYEqhuTHlDNR/gkDG5EMVxYw
M26puUHApYnMg87hLdWa0fDJWQvwH+ruQMB+czpc1H1E205Ki2XMuIal5M0ctTVQ
2BXxNiFymdzTKLd9TUBMXRExSL5XMZNqH4Fnzax3s9p7LEb9YVKNv6Skgrmolbk2
d/o7XL2vJKN5LdepeKrCXjxdiQh6hV5PG+n5sK3XTiWIerVlzHRNhBalp4dlnHRa
P5+i/DQcqwj67Qq0BRiaG5WsHypRuvZQ/tMdem2UOCk/yfWQo7WpVctMHaLxL/km
y6jPhTVC9HfQStiq1zJevFlFzW0BGwPF8AfqfdHskSaoJ6JeMNZ0gwuh7EUWJET1
stJpGptwJsttaeXXWevvE4WapYbHv3KUzWZXbdk21hDQoBo0YgzsfLzHlo7ct+ac
iHIUezf2Hx6hqMuemRpfvrBVA6QMk4oDd7Y4ZquIW7ZIYz9Em88rhz1khP+2jMZZ
/rKHOoyBJdnzbgaFsD4qla/xW2VESooVh8sjGMv2ySDNFSr2BFsvuIHN/wXIXnvc
nDtc3Ts53FdbpbqK6TRT8GdxZDQ9AXlT1PL1oEQfreccBxexHgtFh4kgjFaz/mXr
FA02q4OAAb8/CKWJzf3bn5dthvTa0+yX14y62I8DBkKYFZGgaWak/ClfH2p0x7uV
06lf5xtPbqIEghTLq0G4fcsb8tl+mTs98n2EfzC1IuZsg/G9+2hmy0l7dtpE0w36
MFkUNYukT/VY/vO/VNeKJwi0LUZKp7TGXi+YPvr4aanYB1h98iT5X4Fn5sREi1Sk
fhXNVcDw3TwqYOXRxG93nJAzKTXgj6mxstkjdyFPqaCOtz98dHoc/0wnnrQFplc7
SScgZPAqz10q/nwVQK12wB/sG87tDcaLrolGF7RQui45yDh+Uml0ORHyRumCsd2d
z3+7spD8pNPVykrIeXgvSfZdhKfEW1kC3XqOqbARjEi+dOPNYekf4MH4KncvoRu2
L8UFYJc05zL3qkJiXQ2+htmQGe1kIpMtlFoiJ5KnucsoBNj5Jr6PPzg1axsQnRMT
cewVsNwbm58suY+gcV63N/DiCAulVB/4YLIFWdUun1DNbMSQkzedmVRp2cnQksBb
T3xpVMQYiDvpvU917dXf02yme9lJVKjsGGP5RjVfqjaICByQhpOcGmBCoPd6S63H
5wlG3jeuVIL2v0mVw4P86T8XKoF1HIp33RIg8SkCDg3C7QSBXF0MxsTx93zmACAJ
wCAR7zkxH6yAfGEkiNh3jW1FZko6IMeo1tA2I+Sf9LOsxxT8p8NUHbnOFjQal6df
NutwfH5GCajTCDutrKoD6GWHZ9v4+apOSxFRodyUJE0V8xT5WBpxPWytY4nDmgSr
pUBQwq/i2ejCfa/9QhVDJKO/47meV9jkB2WEMmnpGEG1HXK5T65SnKtwFro7sYKh
0ZosBs8OZWK6pevFVKs91i1Dz3snvuCC3i0FnBr66hanaKuvbdMop4c2SMwrJmP8
dBwb5fcKTkX4mmSXIIa7q5WPPsDPaup4A5xXLPCdLiXEr+FMft4M7S4938tMBg8g
/803/Ti4Fe5pb9vYneVdcRbR3CqgmtWSWZnvctQ/lsjGSWnHpWQLlICMV2gS4OMZ
6oqQDht9a6f79b8P+2x37q2h2RsfA/4LVy3mWbEpg0muNHMaBbAh6VRzmmG0vTkA
XGEBpOHoK/yZ3pAc9R1KeAK7pxCFjcWH9X616/I5YIjgZchPQ4MhfWKt/q2Wm9M7
JnJg0Ofq2SlkkPGia6XnAWUcRZHPrvQQWIYFGkJfoPQ12/Lu/iyvQCotr9gtggVC
vHyfH90PCm41mqDjUcJNWeam+NAbvMWQnVMU/6K/E46Mai79RxtLAIQ8K9xaSo2C
k9+i1zL+pAcSmttfswP8HPWIibx1442GAiGQ/D9rqoLUcFvVaJP/uPxhdyZJRAI+
auDe9grHk7z6Y9AUJmWndk22gkgn1n1c86zb68xCHd6pbosU2LHKjZWTZVcCrZ6N
fCwkEpM3f15bHQHjHZFs31vbEHS1wfNywrlSzpDXs2TDOd8Tnb/8IpQKNBNxOl07
dd/VX1uQPdlkRzCU+Aaw6VKomGyvjnrsnn/iayJ70z0+Xq5LFQuUd8+BH+68Od2N
LE51/kJt3fYn8PTCKPLp0Fz+9u9Y0o/T6UGYjHwyj71sMOHLngyDdnNUf/VA1NNa
RBgdkVCCyx2uput6rFY6BLgHq4HE2gg36k3fcdIYxDb2bnlEmfk7n6scHQ8SzrsD
cRcukkfuxTshNvkR0qIJ99+gkzP0XNaBgkANCGH2+LLpzCteTM692aqcayoJWNQD
79skFSh32vojuRxeKUZDEFomE7NqsjvJe4zv2gJa3aFpddM1DHe8hhsX6ySKb4gq
y85UJ/DN1/1nW1rLsylJ5M5+oShfOXhvNO2c5VutoF0WMRUABiMZf01ryOZxtcAT
4nYvoVSewZSEiHP9B2qTXFxxDJWOv5zpDf0BxKjQCMxN7ZItplGQPQQt50+KHxuJ
PDI1tH1j9VCizG/44wAXt8c83j9aG3rb64pmHEO/LY40lSpvJ702sXsMrHntKvwu
rw0xMuwtqg7328hRStO41FXEpA4wAU5L9+GHpf6PZZhnoSD6jvUM019uBIP727Hi
NtDZ/RilDgyopOtWc3WHGXbYKO+4L1BbgOevrZjjJBW9siM6Ly6L5HIzais22gQ/
r3+jRSSS5awMjR0vJctDVk6QfNh0GppxeYtg3nv58kjQOF/ugC4U3NUdX7bLvHXl
/tptGY8jCroOP/8DvQPsjVX7WkVr3kHc1lfq7WdMqmeLwgoZIHpB/bBAZ6u0x17O
MSJza2R6D2XHVcxXcHPofk8fz5V1g/+FPTfqhdzv578c4GQIwcGQWJoHJ99pQQju
81zD5Ys7cVamYfeQpWq5DwSH8yKRLdf5CxsuAzss0AqUhE8sslEkFOM/hcACDx1L
RZabIAe4GTaguqLGkLreX9BOhShtiWlUI7f3xS+/sPVdgydhbly3AkA1NOH/v30M
qKxb76mA3lqDreF7O939KhsoplAMsR4IFWSo5LSKIYohMpYgYnAIBbF2UjItAQK1
w4YmVf6JQF341uoFBbvrKlKvoq+qdSKC2t4F3a7ruPakhbqlcjow69IlEzPykP0Y
u4YWa7EcF9aWOFm6m8wyyj2dCxUkr/lRruJ7Gzd4sN0xoBxr4XYQHsco54eEKXf5
7PqbAJLX73l54cjolPBb1p3fEMNn9e3DBPbUs9guZ5O+qL67kH9y9btoyYKD33B/
E4ZqjrsabHbMQs49wIykZOSrZkR68MI9eux4O3Roy0AnxA55d0KdAlHIIfSmGfDc
w+QkyyTMLwpX9JGzoYXeiccD8B3WcC769wavQvpj6GS8hZIfp6GmRugklCfXea5A
VN5ZFXsH+70nCrDoRZbawxqfWlT212zfPnPtFyuyxv1XQaAV46ozDbx1tt83ZwRc
SDEftmdXGZVTY5NK/ZNho+XblKa/MbAjTh/qOayQ5JHZqoAVdxJqWyxglXzrALez
M49GSIJu0WYCk+evM/U0UanVF1IyWS/0TGtQ/siv4LM2XRDqjMUjX/KqA8Wy7T+E
apSy5s+XW51QJv/WLo9pUw/gPV9X5L7lix5K6xcxLowQuoCrzKEYKmPl9ttGRX1k
rmKEzlE5aB4wq7t+RbzvDnnSdM2pGTAMntvUqRbE6fey1RCmybf1BN42gUWDAFFG
n4q6Ifp6NGuhrd39kNFXydOyafSx//DD+QVkFwSny0L0NA07oNoDCOzw95LmOD+2
V42j9bgcr6VkcAmQK7+2kiSCU9Pr5eUhl1qBdYnVdMp0u37l/3fZAOkUNhpay49X
/m9rbswyfT5oe74hyQyas2wzGj+UqOEbvRShbu5Ree4fho2FvFBKQlmNrVKIKSB5
j/MFLvf+zfNK3JPJ8qNvjrwJsvJKgdWtMYETsgBH7TE/a0vX2+ITgjIwGNQjkGrU
5Orre5oq6mVJtVrQioYUREhHxi8dD+tmi/oWSBBHYz2M3q9N7hmTqVtF6c3zhvVP
cMvdzpfXC8XSKTTLgstwDnIlfDirqDtJuxDQvcj3EJd8QPQ+4N6uqbgbvQpcParp
BJeXfw8v2eja5D/Z8xECDwkO8qtKHcGJ9AImAZFoqqNhq8tsLW2hnNAvZ6sMpKsJ
sXUjLlCcf9F6V3Dc0TLjKJSwhviwDS525JVzZGTRqBSQ3bRrQXqLx6Cqg7+h4bPu
n2wvNTuLeqkLiTNXxFfHJICMcQaJ4c6L/VNoUrynaVMT/ySsdptLMR/0yxkDZExX
O2UFaoSHI6SUhTle9lsX0tT9SsrpJ8dz77cFYiuY6yJlBj0vqWJNk//AVEHj4De/
oYejTi5uHlJoR6hLPbvfjNXQ1jfZA4PZeh7eHcRIBjPUr7+3eUoticC7+VzIGEo3
LcRTkHs2ewlc0NTzperSbVUvKbT42vHGGB7sRcqMzHdib6N+b7MAFQ4I+yunftV0
uiOZfjw1Ms8G9THl1QApxBVAdK2Shx0tnXnKnz+n3WUfHOdFC+Gl/Bz+L9oLwSS+
FRkciC28JSwqQy0NOpf4WlbOgqI0QH7DaDi7OjhvhKMN/PXbw86PB6dDWFyvKzrl
km6HaTjp49c/XhtH9SzvFp0eky4lLC6DO1NKGDnE9Rv7/q2Ij3srAWrKDJkNdNH7
eGBJiKb+MTfLsk/D9Lh23jc0UCtBEUPHOHETQRt0cE3rvDYX++AnmXXiyrXEZrNG
bD3Ly+f5RP2PL1l3cDDN4tHblVLEmF8fh7E//rTiuArEDV8GLs3FlSw08UpgxHhb
WMg6r2MmTYnwoDzG/4FSTrnp4Bmhru9FZfA3hCitWryevqm/A0NblXAUl7aimv7o
5e+OwEhmz3k/tStQH4rguAucoJoOAFN9ExsRTrBzHbMWok5/riAWwLHx1hf1ypgY
yCEIcBaF3RY3rp1d4Z3ICYCjtP2X/aEimzWsRINu/ZBW3/EyWnF2MM8XBY6vsrtx
Vw/5WWGsUrBN4u4cKDy/f+ZQSdRhzZHeYZV3rTTh97YtCzJUJmCPwCy5Kfy0kUMT
WmgdH8lL57nUEHbFZk0vTSSx9Oa33Ez7MdbmczQLszb3ki1yZEgcoyPKEoXGsd2Q
HjpVyjZg3ICOSNoEhc5E3vXaQksuwn4cPobGyu8n3evR+zUMXK3XbA9G57LnBFBB
ouMJ1EFgGRnGKnEMFf0/3Hj90sdqdQfL5Z0xlOjQsauEmrdwsRNEovUz6Tiaos8R
jnOMOOipGame6DOnHt62hmRKYkdnskd5tMt5Tt02VKWOY/grahyfcQ6DTFusRaV+
FYk7Df9rcSz9OoziFXMsnCOkhN0QatxiEy3vseHV7tA4UvZ1/X71QujyxTtWP+vg
DBrfmbOIpQ0U0grumAsvTyC6qs4zeErM7AI14N0sZ6Oc4NDe7LZhq3OalXjinLRj
Dq2UaOeF+ubEazA/LHx5qZlHEgtzdmWGu4La2OEL3A0fzI4prgESC16r2ZfuuDJE
424DD+sNs4Hatb40OXrb0aUTAXdq7D8lhIXYhaccneikm3Dk9ITTZy1zp96RIff3
ooDfMKYyR3rvop12A+wPS25JlHz/eIb/7rO/+3HY1bxTWmh2Ibk74BIcegv6crNb
LkHtZoNoxhcInmQjPdY5G0cZiKv9FRZ87m3YJNcJeVsfQvJkjIBeYbMSKrUTAanE
2qJyGEdwJ8ZGBgxnfoSukbmaNdoIlAjkLKzP3lCQaCmv1ADdAXlpDMEedOweV70+
YfSwZ8PXsYfDfxbF+aK4a0Nmd30vnOn6PKiEDnbvs2BSYeYCA6AM1xhbZVeJt9Qx
Tg88Tliqth3tZqc97Dq0ltfShnF+6PJIDxxihF2NmSkukDZryTfCWksGvi5l2dcT
QioQkl/1bd+aMg7FccoaXanzHEXg5kz/Hf38sZbj1+VjgnrviOgDhGsZfeK9f4Ax
j5cI2M3PZQuSavTno9HMD8qNMuaYRfaoOPSkqbV7IufDPxkfAP1RhfmHTy3EojH4
1WbuamuHFCo5SZP8JzOF4f6enLvxCLErtr9QaI74wnT/PtKx5j9z9IehiVsQXHgW
cnwxCV7EFyhuTv29ihvfzzscOX7Y57mKlZhXgwzfiAOVM//dGfUWbiiDhFWi6dGf
f40svejtvNfLHCnEw5MIDu8pBlql+IPnD7/rSFsrOfu8SgUQqseZEcS2rnEQ6ptX
BHkZeiHAsj06vp5v9O6nqnG6xp+Bz3bsHjUsSFDO9hn6a7Dg2AewBAGMKHB0mwkB
Iio47/I4vbxr/JnzNy3rVZxcXDiyKomR0k7IeaOQtvN3AQvlV54bgiMBv62nw/Jm
jx/wpIIc8Hd8grJprHzyg3HrpCJtldEoHfv3bJAg//ZpxHXTKm41NU0jYRcrIRHz
Za1v7+RNkmcrr0o6hvkRkYMOHLRO7CjGdLznjBdrc3raWmAuFE9OLU1McAlgzdDl
35Cb0041LEm76vVW6ELOXAUVB89GNqmKT2LWGm2tCzcEty+cPntkT02StWCd2GO5
GgCvACoPMMtXKVexv1uyRlER0sJZXtfynZh7ngK6vwLiTlT6N2UbpA1b+8Ndgf2W
eHANyHc/4T2ihF+opepIsmyM88tgkjmGQSkXQZu5YZU6+ZOUG8Gd+XpqKUfL/F5D
ATirM5rd/nXq11XVfois6ce3F/bznx6LsMzGOWwXKSd2ls9+F7X6WIFsUBYYB2Ap
zA+DF5eYpvRw8j6ZdvjbI5b6FxeMJLwkc45hfDHNxi9rCb57MnizAW/FEc2Vq71m
r7ECjvHHMJD04r7VItpb3/SY7rAOB7+oX/BwFSiWVIgVTOcqe24WVB2WtU6gayKp
gN5pz4X16xhqqSy0j9TugNNg5r355zvbZza4MrdD9R/VGCeRhBRpFs5SobLxvgU2
zMvFQCHYZ30qfDIkAHMTmjGfsCJbo8vWl5vQ97Erq7DgCa6FltLNDsNrBDTbcPlZ
G32HpxJ0btz4V88xb5chOZBjFr0H/ATkaszCAmCoHaBSeDsLHdVlpTZU2KWlF5m4
3OtVbvrGRALwmj/BocmMQQtlN3otOc+imvhy7N16E98wmawHwYT5pWjsxYeardG7
K5x8BFt7GLp9sV7IROdKXQN6ooDiMeM+J5I41/qzJJyb69DBVJVAWgWfU2jzTRwy
Pr4dHyAnybqQikgIfpozvtPZSBeiYXBqRE5hnT0ZOB2pPq002zsrf/tEyPUoaboF
6QsipJLeAopyHdRJIMBWaAIiplaV12lsLGvcf+Q6sgmRXGbHLUl2oN7q5R9HeXAh
Z60dZNyk8rOx24REtDPXVWfbiaucd4Se87QlBitESp/LPnPW8kfMVO+w6hpvXBIo
N+2FEi5kMQoEqlzCdZHL7JKONitMBiWXX6L+Jzij5CanqhYy01XSIApp9cLTNdLV
9N08GNXdO2aYTLSXIJmDnAhXZ0712jqeir9wSHQMfJd4KZkT4WMzef/zq9UsoQkY
S0NLKPGQ9qaRH8vrdMq/plhxm7o58UZNRLNbDvKnpXvD5/JEfTmGiBk8meblVV8M
gnp4dnwrfW8xeq8Dq4ecIwnEnEl5HldDDs+sSMJSSLAYYO6Bsug1azYfSF6aJSYK
J7BCx98i3MiwZpAriD5F8C4y5GPk8zVSdXclZgdgkCUvgioER+NLhZuVj7AlA90Q
GO70WlGzBJuGiZvxCW9S183Z6Oe6Wl3hiVq+vPVQqUS/ACkYIpjw96FtFTAly87D
3j4EBQOzPES1+iH6fbPf1yMLrAW39O9D6JmCQfmjtcdoCk7xdrEFH8xOwB6orXed
WtAYgFZY6qNfVvHnvK340/XZxTrxVorlMjtbhdob1Kzedr4upHyJkr4kTyIPH7nb
eY7l6Vb4kfZSHLupZogD0StHpGDPfXtrcHKhwID1+O9eR/CkTNZQTzGLpDo+BZbH
ygyeaG56kxUeaUPeMLFkfbNF+zoZv2sXjw2g9PhmmbEYJizwDNAbA8meDXgK+hgB
A6kL7S+nLiwPbOfjLU9Iy2mQciFn+2OqSPJIjEjP8Pv6Q8eCdlzGrBVonNq2KO2U
UVrZzcvXlMiaS3K/ZXciMC7Lul3wpmHZhlVjtjOXRXb12z2aCL5Bo5bVMO7NbXIz
C8r8yjynowjCu4a5TrcYRzhoQSoqVUBx/XzOwBiI40kvBIQN32TZI20ZUy1gQJs9
602ImlILqezOkmnsUVoYNvq38sGpKlTlyKnBbkHCnAD/tHhIuWxtIfKCH99loJKf
LCZavwfrg5hsElwd4FThCbHHwRWDbBPUCxG/VAxe/iyLAZYwDhjgMCq/y78Erl3x
f7baqb6gj+uTnXKpLJ3/mC1ePEiCMdUjgFShYKwyk4iUGrDZOqHHOmaMCjjC6KMa
mw+wMmtjd9piJ9ymn5OQYeiozeAwYi5QEDNqsrdRI5PvEZaM5cKES+fdwTZV8CEG
EkyPyLj8x/OafW2GxeVqg/k6w8KPt6OLF/ly05F4Y3Ie8LYnf8dlIIq4tFpZm2LO
Aei8ctMIdfl0Hds7v3bRZ4tPQ6ND962ZoO8gV4lI2nzWiDSu2yYeqggWzDG7qU92
NBZ2Iz3tE1PVEHrMtyacza3ZgxpbzIl+z+rrl/MRR4AhSNCBVOkH/zbKJQJ6TOGe
wUeQlQ6SdlmYau018Y6OyR2A8TIzFsQ0rmEwxNtxvZS97vq6N5gIJGzA+Spgiab4
9k6ZyXmf05ewySrR4BQlBY+Cpht/nkjCnOjRABXwifNWH3cjIZOtwJm/BBAkEy0A
DdJVU9E2iDUbs8yQLRZuwISYrGXGTske3x7o8T/pGA0mME44/SvKkplGW8NUm0Pz
iTgU1vSP4iIPoEG1rg20JPnbkS72rfMGotdb6OTv7PuOvYsqWEqwchjIboHNl95n
UyDmnf7i5nXYKPFZvSQwQHUMFMKoy00p+HwMr8R5Qwf92Rq5w/S6oTvD0xMv5KTg
u08jUukhT7QSkqXK72TUc1WDTlbNSY8hrDXoBp9zMSDKXmVk4Hechvy0iv00S8oe
86K9AO0Y/ZUciiqZ6H13NEiAltGTsoMYvgiKavxu5Gh+C+39Onb3lsLnSRhvG73y
p0VF/Eifslq/3v0aMlqEK6pOc/NWnFqg9OUJhJb5EZWaKOlFPKmcP4CCeVKyFSv7
4nxpYJzOm9M+8jJZGzNY0zeG/d73yeHFYqubA4SRJv6ICE/fHkkzqllrNcqhzsuH
2kXaoPvUI24nruzaiEK6MvgMVx5xeCNhjmD97LymLk2kMt4IDEcfzlkJdRUl5j0Y
OQRJfJMzm0iximfs9H53z2xXGKOPECP7OBsXn7hJ+CkiCHmgPFTz2fsRoySRB7Zx
JV78ZWsJg00Yx0aKsnL4Q1HnMo905Fxfuor543wZC/hj6HxTmzWonPYBfKNk2rMH
aRJHifnEr6f+zhm6zx8xqitgje2G+Jn2s142//95v/i1HuEfh7MoKv5TEnpd/R7I
wFWZ5jPqcZY6xkx53aJdMzbJqJPs2fqgHsOlVW6qP4pDhoob+9KQRHe7vH3Smca9
mx4wioE5lJJj6uCAJgI5/v+bUamhqcBCbSTuRvqzpWQbRX5sbIBf/EA5OPzD+EL1
LK7Q5oNu28R/TJc8e6a8AbYZP19gwbdAy2YPhH8ta7f/tz/fjW7V3mHLryXG1O61
0bH5NTcKi4AFe+xbS1w4WDt05EcLAPKyf8TDN3m1bDL9UiXvFXe0hoIYba9oMlZX
hSGViHvvncHG4QShS4RkrC/d7nvc/FFb8Jar6VQWreujv1o48jteHt4sZeqfQogx
71mc4NmnrGDK0JjzLaTX5KwIiK4uy+X5uFN1fTZBdnWpMCJS7ELK4Xhi+017yRLf
TkO8KOy4CabDlTAyYKS6VfhGz3ix1APDuXZp6u6JOERIZavP6pKtnYN+wy207CK8
IxYWHkEfcsYJrKBNKrY+hGyS8GAAKyISA2QdOjWgMMW7CiOD6cZnLyrofyEGsbV1
hbk21HWsuQT+zcsXrjBQWjemCz3cGwErgCO27BFV1R7buGpXcJRISMVBA8xKC19T
1kNo8/JKjVNb5pYRI7zGRj7bmTlwwBdgTbVM7r9ScaNadgi5VtC+BtEzLjIhZtxW
ujOqOp5H+t1P1FKCDyPsF1WD9arud+6XNHN31b2xVZ0Jo1cFYP+Dj0FgXD2/9Ni/
U7gjgsLs5rYaRABE9Xgh9zL70YnonOrYQQ1VkMNdG4yYVJBLng2z9Th1gx/VRwhm
sexTSRtnp1NzhO5Xwb4X9pMxZvMlsKNgDUJjgbpcL3yRLuBlhuptHHgH8ReZeve2
PW2v2kjWdY4vUrrZdi2S80L7sv7CWzFEvYB4T/t8eFxcUH5Yujh+UKkGsvMHxA3M
N08Y6axvhpWZ3kIsELccg2IZ+sAU0ZRjyQAFywPEy96ukht3JkjYgJeN/fLRM8Ao
rjDl5zP2rc+5EaHD/YUUKL444pD3OFJGgYYAR/ieWYsILQoyPpgyNIcDwoH+/nWt
A9TrTDSbJVtS9ha7BAh4Y5KT0ceOx024PPa2bYpx7naoF7zhTCH0cOxYnB7xO2Ci
22pnHhRF1qWZmvnhlZr1wPPIoGjlKbpmn8WV6PGSxdhdLpeGVUP3gyU4ZIgJ9cGf
+epJOJAGtTlouwCyQBiO53PHotfXKrv6MjioHRc4rTfRo0iieIA6XIS6o4mz2ovc
u5zJAwWmDXgO3TxsKStQrqUcxLlXmMgf79YlBIGKAjrMH8q4voidwRFPzPnYL7C9
Xlhf0mIyJd1NEb7XuD6zs08iIr73xkAHJlsznaXuhgFu/x/9oKJjuLipSOw62bE8
nA8uz14jPSAN3yun679mzgmjRXrJw1RGueR3D/Col89eLFbcFAv3en2IFGhr5COm
wf3+t1F9QYtHzaMJvVuTwJi0i/7BQtQDwSjgMoZ0yPLPJHuqY7DUksbudTwJPaUF
0B0wbaj9PQgWt8OqzW5cXBvqDigp80WFzXeWJ2fS8UpGsswQqP8mdKRa+SSJklys
Nd4Dyzjq57tcN8dpw+WOielt6RfJyllzUDSBQZ7lWMOumieZeYATe/4tUozqaQd1
Gw33rDtWfpbHr3jllHdUjB3zzG+nlZ1W5etl+8FX+HEqONWO9rwyGdGz6SU/8K5s
ijI3vezMIlfLDp4NzWBZ792SvIiZPY3vgZh9mpWY/Acx10nSWbQ9+eKfGZhNaDJD
1UaPz7YHLOZNXT1uojllSK/OeFpupHsKj/11W2lblNmpQwfCTG3XRscMZkaHpKqY
gbeJxxBkOyYPfOKTwyavOX8KbFvzgj+Qm7jCJXibYJdy/Kxz/gbxkHW5K3mr7fq3
iwIqx5MTegRiK1cAD+AZ+VwdiTTf8x08hax42+Xx0DWalTSIeFzYm+Igj3a5H2xa
Y3+3jScThpibg0Y74eZrcLfZfbxfFc7dpVM6evnExlaIWrs0LEydjmbQ8fzhP5wK
xzh69ypGXPtpB/muqyImYZBTXi+icy54Wk+lfXNPw5Zrh23BwaRCuX2zmQAwrvru
b0QdpIE7754F96+acD5wf1kwUeOISktaABDJlCQT3Eqat7fdR+NWWAgIq3A3Pof3
qenAopqUUrq6QYrYNBMF4ILYxwsqisO7cGHGKUuhjo43cKmbUoyMnbZHazAG8jxy
Xr3d1EqZLJjIGeN7DwG6FMSRlYbHTDtw7Ag7dND+3QEqqXIXwZ7TGOzPkYUYrNzc
QH/DIdKlH0+6JCxgoEp4p0vOrRruiR3l+91IhjX4mHHNfr0amLbNEh2ByLar9pDt
n610feYeT2SoDxEC8X+NBl+TKm28HXsOFsoi7GMMOj5eeZyrTWJO9dt71tA/9pA9
SWqIqVoQcNyscmwCdfcrV2W9fdwHtujhB7sLlcotawXPTAW3mq9Ngfx52BfdcdF5
t6r21pNphAlAeKs/fq84FHeHA2ellMNdAWKO0EDomxJMgfb2wHq2nbg+zJmwPxdl
s/em9cqIvOXC6kJPM0vtGKHOH2gsWKyq/GZ6CtMfz3BvUu9LnAEyWmCe72zUG2Cp
DeXaAL3EFO07KYPx9vjrBwlpcjkF9EiPE7JA5SEflnOiYmTVr5XUz5b+GgVluBd8
uuqlOV38svGbsALcKV6xp7QNrEk+KtHDdoQknzkv8rZdfjOOfcYZv+2/JaHLfQob
2pVcD37I6XQEVezQJgbMDk+PFzqvEaT18mXucahARf+mTUi83SMzyLVMqyvOVqI6
2UEucz6JGdOzfr4iF1UaqxpZ5qge+1p+s0wMrXCPUUz/3Er6LGIUhPpRd94hdWvC
w6enXLn7VA5hZYbPFVvSl04f4vQFYSLT8oZiOL8AG4dTtieDw4Rk7xlgZg7iJmQF
wbR6HetSDkjTtEqrQt/LWEToTAUnJtih+ntPuXfOAZ9jIw8Bxc/v30cGgqn+4NeO
lzMuZbrUiAmGwsurtqEzUuJN8KFN0FqdiYlNHP88uGLOUZNxPqzApRlwnz4L/BJ+
7UHDNt+7DRjRZavewEONyCkQ6FrDcpE3n5icfqHxkT/afKOYHPTL1kaj6fk+x/gP
rB5QANdFJGvY4U9L/MeH98XnbV64NhKZu/x7s+Wwy1e+oYeKTgvejue1ocziSQQI
tkFVUjQIJ4GjJarIcCOqdL5X/B/zNdVkz87gWvADREUAOXWGLHzHXCq0TLPeau7F
h7xQMw6FRZYn0LKoiN7LREHquDeL0zEXLn2JVTsFfYnYMWA4XeawFqFfE0osd68S
PtllioIbYBh34/2ht/Wq5KxXJ5FOx+Vu5gaofxe79mev1+T9Hnb9YEwI6KrN1UTf
BeTlXAuzkag/xdL4p9wHWlKELwc2g4AGDwMJ6o1swgEhu4fdGajTfPjQekNdfexa
QND05cfzXFA/Y9ZvfrMvEm6uQZlynGZe3dVdmP8nDpAqCQZsz5cqfe7oPSxB7V6E
d29PRrlRZp7d96WOQWhUFf19nAoxmwM8p49iamsJR1rwly+rd0nFcXlCOtZpVFEf
rB/QwQUBPaQpjvop/jcj3ZVDHDc5S/2E4qYnGp2tOwBmGiQN2y0KzcZQN3MceGSE
1KszshPbYkK1Wr8wA2AbwZvktC2KocTDhb/clStR4i+icODOuHlK9BjYr4CwEGQ2
MLWlr7+NS5tZ7GhyNLxUJRm7/653CohhGz0hBF0Xivj2jTgZDKHWcVTeN4YBrCU+
N7W21Ann/uusW8tG52Df4yAJfAz1XupqILgguQEpoL+axvojkN+e4fpWt3RM/YCX
Dd/DlD0IdQCYVP/vx5mRbbIm2TQ1th5zAaPUQzy5yMO6Wv7R5blQmJ3GO6ynuXCI
ZwXofpZaawdN38OUpnAP6IZk3CPaRTPf2Xdyny/W3WnXE5//AhBnV8hXRZ7/I+Ah
vg3ZGx5oR5DaiIy7OxxBcgjBClthbHxzpNj10n1gVELVKb5+2yhArLAd4oldhyuF
+q4F5kARpnhGxnmyethwU2BvToJA1DrUvuDj0FGTC/MQfcsuzZ3K1TaiZctSe8pT
Jw3ad5I26ql/Z+JWemUav5xF2fuCk2qTThKvAP0m4s82DohIJ9k2dRYD8orOKnZy
+EkntTGZ+IkepYVgStHOGnfFbA5tnU7OYsPmglR0L6JSZ5OaBUCVXJEfPn63/m/E
6PwYbrN37XCi2GY+pKE88uDMKQ9pAmR5nhOopcwESo1ZxGbAOy2X8f2yGy5IXtcF
+I+9fWh1iblHdXSRlBe5Lm7u2Wu/Nso+jl6jSEU1n8uQkOVqx8V0ux4Dealq03Yh
D0Wog1RDg6XNGgXfMw9td8iLY+fXfKxmxo7l+T97+miVqyykCYmC71UfoVxd2ZxO
+EYTJLNhJqFncQJ4E14F2KHJ70GtFCAOL8nnHDtdXcdeqNoqVCGH23txLo2llT0v
oZ3Od1qyvQwm05Si5vVxHqHsPG+Dbzz3iAEewAhltCukz5DHkHFwpDMBUu0hhXDC
V/QRAmuKwaZINzYrem8Rv6kWWfkFPI0l276jLcmYsVMy+tL2SWnrjv/tSWG9vbHB
7jXRXX+Rf4lXynBnJQMiorhMrbiDkzGLP/Ayoca1gZPkYxS2YWiU1lEJWLVwxw/3
10fnzmzqRLgNqSGZRZKnIVbE0jbOo7aBaFcqwysYjwnyDq6c8EuHBUtv+tKuVR5Z
pLetPY86g+q2nCjiPBgQBbPjm5VlXAFibzUrduBiAgChlC1WS0NUVwH1IEZ785nb
/W0iUPqUYnDgF8lnXQfAsVU0DGv3Ua6Q1umSaaKPhfe4xl+WEuzR4R5LQeT0/Oh6
t0drTtWPiNPgryHAQ/iUnT0lFIhQpnCkg7VeSRsMd9/gFvBdoxssHKofhSNvz9zR
4yY6WnnzMvnP6cxS7jqd2RfSXmmRuOr/dYYz03L7erdZfxnmzSZ8MSii1t5HPK+q
Lms47TPiNQqfMSttbVfcWr0psnPHvu3ewsJJFoTZn1GWGPw4nj/CvUevC7c+O2q6
q7A9bWvCSyunuiwTg1t2Q82ahZGpBHi3Jjlmj4MJCKX5Ts7lAm8gl3oXMEGhLK/u
62fkAk3IQnHOD7KxijwaOmD3UI63qeY1L+quz6pcb98M3PYJn6S3VjbfO/ddBPNc
hmZo0nl78hxKGuTJaxyvFXCJ8QKXgaD9BHJua7xS8TvfR6irvup0XLdstHnYsN2h
LTEVXUU1bPjVEeeBOpG1SYfz0o0nKrEYesYa7fY5TVHSYJ4KK7XnWFWXPi+rNwSb
0EYF0WWkA4SSus+oq+vw7swypyu71zUHSrkSHjgaeBFeacVhgWULWf4mkynhCXL3
xcsPmCTirx3EXVOW3b1gGcPXRFsi22BoDIZ1qp8YqU9niVe+Z0I/Dt23lwZf7Lfj
2pnxVaVnYXor2wNbZoq0dR4PpRtXARvTL9k1zok9XElcpZ4x5BIom18yxUJKqI+/
Kb2t23xuBpEAeCJFB33c/cWt+jOb4vkzb0+QIC/mABtkpQraTjazpB6UiEJR8vBc
h2n4GujhFmpKpdMwc6YAgG/6kGVs6c1EwverKwRNQzWoUZFt+IaHWxh+8VlF4HBB
DmdF54YjFNe6PFE4tYLCsvW1qvcOh7kHwBeEVaWxF4TSJnh2wlegsTqnpdhx5tlm
1eIh4+DB+3YQdwtpWLHNXzUPoCp70Ppw3Gung31WHboM3LV79SuCuiHRTMf8GJ4g
MNh59TjlIP1WvUM27LTe/iEOtkjbSqnSb2ooUMKEeMK9KNGdtDIckst2O9rt/jmL
JBd3XRf4EObGBLKAr1b6wb9DWAkGc+URGlD0VCQqzaz7psEiqs5lBqT1XjWX41T3
jAnMiN2aMp9ApsARX+zeQMBNk4qlefqyHJmze5l2VmUGmDYZEyDzAkb52VKUjQEz
kHlmT8b0HHM+bTDEdsP9nJAThA5jWVIU39M5rniV75cciYc8xHBgfxonv1vGRtl6
/Fa7ZEy5T4Jcn6cxsypfWpEQkLbGxIW1qKF68mtcju5OYBCYMNWscANYl3uKL/0A
Qq6wjP0ZmjZUehajq0QFZahQavYmEUQkDYnSG27g9dSpW7uq42HMXy1g6ps+ktnt
o9aM2BDK36EQXHmkCLFW1s0n2tezY8UPmcxQnNG52WSWM12qFnXz25+mbTDmxFab
fMe5crb8cwFZCzklmTb+1Fotof4FQk9vWCzvRiHoWcayNV8sAkekVdCSp/Vpe/ZZ
ChU0o3XhAnclNBcx9Tzftjt+9k/TV0DvHLIVNssENyPa41sr8Lwb8VITGwBadhAD
ZNUNKOFIW+xaMklCYaSEqAijh7+IX2ofP0IB3F4QW8g2ciKxa34RIuH8NsOlc7W5
zn3O0Hdi8BBARWFeOvkEXvymWhq3oo48vNkhlU5OnKX7v6ojnAe5K9dYLOkDv5U/
y9AMpMv1AjZDjmrEiIPviS7VyAveFik3xMduY85vftycQs3R5Y4tFgQyRahoN6Dt
EMm72AozJu2RasknksmDKuTao7TIVNfoDjEJN3Qj++Q=
//pragma protect end_data_block
//pragma protect digest_block
pg4Yk+ZZTXiffHheB3cN84HNRSE=
//pragma protect end_digest_block
//pragma protect end_protected
