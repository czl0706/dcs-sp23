//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/IVXrwq+VGILBFy3sZ6sO5w7VM4eR9ej2zLKWHJLZcSC+xmJnnHTqJhFnLSWoHQ8
63MCk9P5xsLdhth3h20Tvr1KUlfXrEw3y6+g/a6F5SAgwu6u8OsBfMZpB3tnl95f
FVxjEK45p1SX8QIuMp3P+jVQxGdbqnt/maNbBj8COWknSAElDlhZIQ==
//pragma protect end_key_block
//pragma protect digest_block
7ZwdU3R+n+DFDw6ofd+wsfC8WXs=
//pragma protect end_digest_block
//pragma protect data_block
gVNbSalXOX5nsgViqU6fW6zBjEiW2Xqo71ox9TSbeFHvkem9NsRLwqq6mhDXx7hO
47z9v2aQneNR5z91BOD3N3K3HcvaPOe5HB7zqxffT8Jhx1DNCjoY3rtRwxcr77XJ
rHdO77KvsPlaqhEmmBuZY8r3RQ2HxopRJwMT2s621JJgUeK1vl/9xVhwPjpQ3LSR
pE9oy2oCG5/7whERAV1CV8JuLj+1UeqVPhJZ29FLOG/J9Jw5SGi64utH7f85pO/O
Kg//we3Pohp2IfnC1FT6M6EKO6MyqJI0EG6R8bnV3izEZxPTlDDu/W6AOqhg0VDb
oOl9Dfiqke9Kg4GEGU1xiZ7MSVOIweP95BS81G/djeywL2EnR/am/6v7vZ6l8DSK
kRql2Z9IhVZoTWdrM5RfcGVINFS7la5SGx2aQEK8yM2HNSM8y+e9AmYmwHQGTv/z
z/5GujD3nNmkqjie/b24ZCDoFrdD+l1uUJ7udqmreG63WdDl+K6F5ybaYIj97fju
l/Hkso/lQSsrSuct+mdhZU/UDOL/OBg+qe5KVZE/Q1ts6xwYpozLH0YMisYNHx7a
mk2Z9wS/ohiyCrShkzfez2qHcjiU6vuJaMEVYs/84gSskVTEmsNDotI6TNUdhclm
3+ThcE2KomWiyNNfEODW+v/W/Owag+3ejlJIOQgCmuMw/+TEOqSsxeuPLb9lk9PP
3MPl/j/62i/RQOfxGxyLLm2YCUUIpQKsf2cizl84HSNzLgCrZ7U6i2IqijTV1N3n
tp3SD4EmaYLoFZdOkLDg1u9AIF7A5Flf1nM1W7y2wb5XF/EDrsIlm9Md0fiQkW5k
23qCBmnHJ1Y/9mybPP/syTd4JM88bY2ZBaFwODZwJmTTOf/9PRCtBPx+dF0kbYE9
xmTvg0LVd55ykDY8W5lTuvmRc27scz3rLUF0WDS4ES3fLW6CHxTZ0MUPJs+qI1f3
58h0fp6O29PkVL474tA/5/Nv978NuPOxHhnloYxXuyN4L02ficUiPlQtkRIFb9ZY
VH374baNxEfWQMvZzzkfVmZrtroxVRNh+SJNIxrcTXsDN2pelg+Zn6X16TTEUNVY
iZdpqh6ddPxZIgrJKbYFdvjYwi2wp9utzXZZgBvsBCW6zWNuniVowu6x5XHXL3TW
yeBlY1DeieMOHuqpHP0b5PS8tyodBjLctRN5W8RCQEswXjq4129gQG4Q4a/I6+Xw
tHoerwgyuzLy/HOba3Bk2Vbb9EK0ugeuO0DvF9Ty+6R6xwtn+bf08MsffdMQSZql
8zdBYmS6EPDtr0W7Oh2Oe85Y62Pzpn3kHNkm6UuP5f4Y9kZEklosJdEgovCLMulk
Or2HsUBNWBO5saZfn6a16bErCMPyd2MUZfU/zPedwPUZqzLUUICnm5eD5q9r1p5P
c/adVZnIq1b/o05T2QctKhNwxVhTMJYaxWtc4W1X34GYpDpd2oZjzd3mRQ7PXG1Z
r0NAk68A4CtoAPnuaB4aDUUhl2oYIMFFRQlndNUVcOYdWGUoKO9RRjL5I8zFyP3q
OQ+2uN9E25TdINKjgMP+ZfUtdLW4RQykh9bvoYG/9XEPR8p38AP3tMXVZFHJKs3Y
o0xNPwpi3nKngSUSo3F9avAWhVcpV1g1csTi4pYkEuscLIhnQ8NrVeIaKKvGKrvY
7CLWRsI943jXUso2bXeu4set6jJi8rTYbgkJM1g164oZM1P95P9kdhtCTVmdoEK4
VvcEzX78INE8xBhVpOcJ/Lh+RwNvSUd/DBVm/JkQ+vaa/+9xv4DqaQzSsMWzc7QZ
+bm2FU25LiZKTLMAWQ4uqxNV4dOOf710AGd5x8Jr6B7DtsEO2sr34YkBsEJw9aUF
lhS4p1VmfKi5klVUM/XX846NK9R58hkPHklGWdkcyHge65DsW/gxrOgG484lo7Gx
EOFGYtIjiWNADDMBXcwHg5G3EGHkSnPgpAALx0bgsClfvSkTJ+K4mNXoFqH7bPFK
HFkmbyaMhdzl23qXiYMwkweMpDFLvBeVte+lABGlqyhvrxPSGR6UOSRG+b2hO4k1
gvI9VqsK9gYzZw6UxXVbWFL9oE+1JruRNOa6yqIkrquPjHMV/u0UwDSG4ef39BLF
QQtllMP3L6VnfqBpax9VLbSfKnyOOTXDbf4TE5rA5wSDbF+KtHrvGEwBPXrBgEyn
Kyx8ss2Vm6TXjIjcnjy/WSDDRfn3txRWv+OU7ZadQqTKOJI0ka8n4raUJGJyW0NH
GLS21VEuRZWUyVh+LFcDQ7ZtP5obX4Ja8zk1buJvrRzWKpuHpi4O6OOyzgr6jWWe
SdBADB7mQ/A3rfKZlfyXtaAzHb8FVzAaQnh7ycrpAN0szmg2nbRPAFaThU0sufVv
KUfBgjrQaDEeOOPBmjQShEqESrhGMmnff6a7jJk7zF4ByGSdS2LY1rgM4QEkhj3l
xK7c4q8RWCrrMN2vq2tcceQ166BDLf3SHVgnXbZJ3fD9w0RmkuTf2WVaZkNZ7USp
i+HOeOLrEhf21E4oTz9pn8fBr2/ICx4aGfEc1RvU2QJRDNiUTnb34SYYyQCB2BA2
oR7fpS9a7SIgTGuj4x+BH8Yc/hlIlUjfpx4mDtVDd6xL/J+aBGN60ZYsW0Y7Mj/k
U1gleouRW9IWN7fcumOoF2R+x1sPRtyLjxdJX+dCY6INvM313FAz3dw2aoY35XP8
fDmIxx23m3eKJVi6PVGxUZyKnB11shrf25kK6Cd+q8W4CGiVQZztxHPXHB+kRS5e
Qbpf/5bSfy/dR5jComjqWUApOUh9noBKq7ucgT/AtfnXC1GYDKpXMXe3lBpwkVUf
nTZA/h7vnOFQeV9EQWqZ2wFIOVoax39Eh3mihQN1S1QLTLgrkc0B5uPEhcxrjWES
1n2iqpg6Wyo6hnwvi1cRvu0MJDi3bMmCHCcm+wijLNN1pm9CG/ez/EluGHFPNqX8
1+7GtXedGqDZLs5xsuXYIBrU8LCoTHsKImJKkuR1GReH0chkBxxnHaFTeHOyTBjs
G5pbu8vwOpYvzboXDc5Il2i044o/TPt+b2oH5fyfYL2u0Qrn/esC69VdCMRY9UZj
A/dlI0Cvm1GcdqotT/hD9iqeSgG8q1w35zKbtwKuh081kRACeNLYa6nB+3JtR6Oc
ExB79XuhNRanpBtWCTOh3wj+lnhHqGp/wGzpshUjPnrcbA7o7awAQnTpGmga6CLK
9z9K1YzcChwTVPlNrk/h7Gjtyppzf2O07sS0IpBMHHgPu89QmQsbNh2QcLosnpHu
0hSkSz32BvZF0REqZ7kcK4LTgYu/RhjXb2B8sg6VtY6Qs6RsaUljJtbYnzlLR5PJ
4Dsp9pLws0X4anZJIByMFs8x8184w7hrnv7mbk7+a0Kai40gzyfESUvsSiB9wKSY
j2VRuSkI+JI8CRlXCj49uqTMJY1/Oo5kZfphDR7ehrkO9VtGDHrbtx6dat46dOJX
AcFAYfqEqYOOeiQOJZ0G9anYky0ELLErv9M4zHZJ6LHPIwSlpdhOomzTP36ujItR
PwP5KWUICNV/xJXxrviZfpOoaaaPpE2bT/auD/L/WD6deyIaWcuERgU3JhXqAa8s
R7dGaekNv7wMVcER5D1OzWwkplSiEyWHby5BguLJ6lgkU0gE5S/Ep2T78ZpDUBFI
wJh1jLPhkGv1BkgQq3zPgToSYh7V81dOsInqIRpqFJYTASmtrxNjvtRVfxcB7Lwq
E2mlnu1dTApx9GGovTbiDpzGT2MKgjYZpLKmRg/Uixdq0HseES7nFVGQLxqrJ1Wd
h5CBzFj1i59DFUJIYuAFHN5sL3Sadm6eNriw2XWMRHadmtzsU1785EEylTvruRPI
ZoL+hr09XXCabe+3vkOT7y+uv55trk65VreB12gNaeYz70Q7N3m0eeGvW4VqupUc
o/uj4pJUNjIasZ9sOCzap9Vczk5I+jlms5t3WygdXaCsV9XrLa+qC/wPOwaddzNq
Q+GUz/ZAfIo9f+YRl4uFPavPP6YR5iCmvDwwyplkZThhH4a1dfrhgB9MctYga6yL
6VkGLMtUf79xGXcsc5pb8CQr7PDqyP9mzeCuO8AC6OTp+ZZEy2E3LvGuBJInWXyv
Dt24d2Ecm/ryp1J2Hcfpy/n3o5hY5a8A/IFIhF8r2kgfv9ICk+MaWd100GO9UFb2
Ja+A9q29ANakFO3ZHJSu8pb4Is1xhlpKqFmEIavWefLNbvMfnX7mIurYIvrJ+lA5
P4/ZpwpqWLYuLVXnF2oRqLz6sM8Ki5DExPxgpM3MX3Dmyf9ZenzgVuD6HWq/ewrJ
kFOwK+IDSVkIj3mcTXZiRBQrnckqd9CuQrHfCSWccHL472S/pOtHiW7fYxnvtHgq
fU1VG9Wx9T9/rFXN8HFxjH9m2l9wI9N8fQPaxuSTdUl4Yo24PeuEIA3TBshCuZlp
6p495VdEoqbJc2yI54rrlEhxGBQww0lv8DGr4TCtDopaNIxSIE+Xd1gVQtCylSLr
qYPYCtzZK2XeayHy1Ke28gFr+9tmPufxCEx97ccHIiPbZ36AgPPqks+FIZ15A49a
HebjVf1f5Aj82Q/lxxMitVXyDOWcab8S5eZY9/S3WoMhQqGz1KPGDyjA4ioBKAOM
1nH0ltRDH1GxqN8nO/rftyS8yp7Z2jn0TQ/UyTGISgDa05+9FE5FvfB8e1T0phCv
gEMrVCYujPh20ySdXjdB1tfU6LmNMPxijVxzwqDV/yGASnTzzEGkaxAcott/JWuG
tvCItfOAo+J4arPaPKFuUc43UqVsmTuXLQEmcX9DpIvwM92lv7zifg9hNPvLe5iE
0XM7OCl7gs04uMwI1D7Pyo+WzlHipjZ4tb9ny6hCxX1tvDLDYEL2NWODcC/e+GPt
9Cy4RKLtDjUJnxvyjHZbE7iGAaNcKU22uiUSM7EvZP34xAAHwEgxye8fG2CcpZqh
z1vEb+oQDfDP1V2B/0mQaSINoIB5PiryKrxaLAmw3Tz0ZWQzhN7cIHlQV8Wwrflx
icIm/e/zLV4onFi/YXee9iDOR5TxTe26y0YZhzSn9ql0LaZWOxiQ2usF19I/tC80
xXoQjRtsTerwiKjA/jUT3DatsL+h9AMJN6SEvSyDoT8k8ycAaZIiJV2d/HjAKPtw
HH+JbcegKWYqaxNQncyIxk0oSIrN6DrAryMb1Wr7NshMhU4SYZADat5iz9uIrZE4
FI1PxdBfCt+3eNnUwTeofujhJyY96F/MdCKXzGqr7vRFTm1duwc/bl51UXDNjOah
1fe3Gmu4TCwUYXhquoZvGi5PXXF/mmVBQ/xJC6MYGS7p9WjSiD6CnPOA2wSm4rpl
SzubzyTP1i+VplP/yM8+03VXm5WXaLT/xJfogmuDpopKqtuNxxewCoxFmjkR6BnE
f39DVLJ3JoS0+M6Ac08zP2GRplFhBlrPlKipy5S+3K2LASol8G/8gtg7rhCmRAlg
UkJlGEyFYLrOiRUVTxruSyeGubFfFhBrt2RnTnAFvfzVMGercNJaiDgfnMydjvye
D8xlsS57JrwQD9cPwywwxo2e8kfj7pjqTgJJF/Od7bYSN7eUDTbE03tgYoBXSO1U
aONrCzXWNIPDlPm3+Z9ykfMxuBEN+9Vuob6WmCsUzGiNfdFLRDeQkltrhrMXqnPS
FMoxvGvmca+0I6bcaCqZDoaIDPaORvtgqnzVBDUucTDtOWAFTxp7VNDSzb+RIqFc
dt/0V0vniO8ATgzt8MGbc8avmr0ZToHxT4pYZuXQvLdaHehTwzddkhXtB3VcJbjR
PqL5jWKD1Ldj/jwrlihf7idkkr2obqNuxgyOKYFTvqvuy03Av1np0xkBn8Dcl5a0
ACKXt+9h92K4T9WzC/7UrActA76W1sWjnfchmCuhyBwSwe4iDiRklS0S9LHzoRhH
+mAq9XI35jSDwKGu2HDvldm3Dv0gMtONKjz5d70qozPfayvuLTbTrGtPfZfxDH31
dA8KB44degDaxbV5I7DUER8wry3BwY6m00OfMQGHdgFyS5C+Q/2bO5RZwLI7nB15
bF42Ok6CYeHvq9gR8OrCCnccTawTfo1AfmQRiZ4iaqg5DXXEOQ+9+HnKcRnD8OPN
9RwcTe77k+bd3ufd0SJ6dAP44wcrH+sVVgDZ3A1mdbaNrYUyKNw+a1di6bYsm4Ln
qFhY0sS9XygdRHzcivwT3L7B7Bh4KnsA2vtWvKDyjcytD1TZlI3HZX8IrdmPiu7T
8iQZ40c56OYHQYpd/os9daZs6VWIafFuipOEwumtFbnrpXRRJ8ndIrqa47MsN2kX
KSf4FXcI2rJ5yhF5JIgSN3GueO0CKE6CSKxft2YoIhGp6PFE5QXgv8vyyLBkCLCT
eA6CMm+3JR6HnzG6UtwnDhbPaxS/YgjHDF5jbzIdjV800z820ra0yyWqEk6drb0I
czD/QpBoS+AOXqiwf2R9u+24Ri4/pjGXmC8WoCKochgrpXg4o3AYRKTlqrZwo5jI
r1sxXBBj2gDGBJON+S8WWnLXxyAPR6Pgh74qniBLhWX9lBf5/H8jktfxVPiXxalL
9M9aPx3d2vi4EZfR/0moJzovIhChrDsILzgl7t+hnBekE9HQJp9Hg+kVljo7F58j
QtS2tS7EIN6Id/ra4jsyT7l0/inmmlxNb8X27yUzeG9iSBhdrOCaSAggxXqw6I+i
qMdKtOwlrogyeCDTbLaEb6LAsTvUOXyq58CrxxLJXKO7FSli9jPUdBVVcfwSWEI4
WQdYoKDyx6yzZK3Yuzr8D6Ct77yqiViy0Cw+O0IFlNE6R1VivGp64QJ7Iq0zpNh0
/sjfVu8sMj5F8SeOXp+1BcadQgqG/HnoPwQLlbHXOR0ZWA20zNgiUP4/0uD0qcAj
ImMXoKG3R1ETClneRiEfvHFmWiw1aPoItexeg78+AdsltvgKW7Wb26EGwblD0+66
cDHeWSLh2mN5LvmZDnvgTkETaUnPsUO9kCu2j2k/LP9umPrrOj6lrj7J+owEqiLD
p4FBpnVsLKW5/FeXqU39r3LzOpVJFrkBt55NSyICjojDPjRrq4iSASkmm2D8KQH7
icRQngCIM5qlOgn4ymxv4KhFjcVhD+JwIlLGhlBlTOOoCkC9Puo1KiU/HOnmfvhx
NZDqAz8jIUyduWyS+1Ey2J3QaI5ehQqROYN2SKP1oyQthqAyYCpqG1a3pFOIN3D/
xTt4in7jo1DNXvHWEC8Icqi4EzE5jhiAKMPAXh1RfdU7XC5Xc7/T2tPcGixD/4r9
GUzd96K7QSe4O7bRFLLf2bMQaVH45qpI5LvEHn0xgh3r8C+JVqXU9ahOWc9ZjurL
Las78ZVNasjsCfPxn7pc71Ns1tdV0lSGO0/KPtobeN/31TiT6GT3ER7M8s777vhs
mkfWvM6rX+6WeeB5CtrWiIgwrmX6HrALd9/Y/cbVWdffbmnL7edfRkvFsoxleh2q
1s6Xyd8lF5/AAGqt7F54McZENZ0kIU/bO/x3zg0cUBvWVDkdOpzNU1ujDfJUmhJk
bKLeiQtQOui6eE5UPUMs58qVbPZgtaN2avEZQbG6ULphQ9/ooWEJdnwNrOBD0xaC
dzfxKYW9WtTxcg1ELY/59zlRRny4X8ksbeyj96TxxsQOMQBAegyVHUcJ0lFWz1DS
j0i1cIul4Uc4TwV108tsITv/jMF+8tDEW65j9eB9MkzsnbjrFS0lMY1M8+VHgztW
jWGMDLywiDuLFp2I48tJ8XUiWInydnb5oqyfo8S+He17B0EBClHfYgppwZ+qWd48
+YEISgo40xRnhRiuBxP6rb+tem2x+EpL0D+5SEiaOnZjRkTjVobcxsmeL6+3+Jc+
VlhS27TedJMXFq5p+ISGycdoJn7razYjT6cC0JZRgOTP5hz9ULZevxsg0cEkz71d
JrmBwEgKTmZixSI7XBYKm3VRFd4nHqDq7bfeE9oPzW6HT1H3uUs5zl73fZXwSiMt
BZxPSU1owB+mtFKP7xL0EyVlmWeOsLgpSfDIGwS3PgpJ2mL3pd5zNHNsoqIAZ2TB
I5k5v187TkJ6hK9Zr/EyUKlD0koEsVBSxFD4VGbttOV5oqSwoqrj4DRuDc75zfdA
5uqmANpotDt1Z//jsppuaBkmna11umuXs9f3EET2NmJB3hF2JgCWB+K/+lr8vGrC
eZ7tgBwcxP02CAOIGhuiNvcJNXHYoPjJyTbUd/G0/p6RVVeunmLuO3nk1S78Fw7K
G9gX9ohFg3EeebuN5Hsow12Axoe7jS0gwK6mxeJrdgaX4M0iRQkohkIX/vTXD0Mn
FvPwmxrChDLULsRXVhiqp5k+0zFD+wajBCpTDoH13ok3o8N4O6NHqztjhQaYTLZm
guC3JPJJyAQTI47368Zfv5dl/rkGkyZXMdHXK8leodqPhWTnjqgxiiazgscu4K8U
ruQ9EToWRB6gl/xml4ge5Xgjv9CbJxP05PPZGqTlEGQLND4ErYf0mCbEgGti4n3O
yWaMFi2o7DrukBNmhfVruVd0dCMx+T6PpM+8hsTTWO0uuC1trYGMqUCqpeE9GmgL
rgWPr7p/z7xK54vJvrgITLv+sSjb8He3JAqYahKoyOhQfvra+gIoFtV+bMc2mU8Q
k+JaVevNuFRNBSjRAQ+PbT4taiz7XGSxNkbkH6s84DUdbMJTaj8ltpdSyjijNJIv
hvKGNRVqg1Qa60TJozNGdNQ9xEJi5xGqrmgHsGLyETPNSIy53LtRAvUVrnhS/TcU
L8ZMGp9GLq9VtTA/Wi/udsA6l3LDCJ9qGk3OU/eIZ3wDA8Y+OQPYbmYnIwgVNaAf
rmFYhJXpSIrTO00y8U95CfESwwO9zRYKZxTWEcri6REPH4iOo0H2n962eIf4T+7o
6/EJzAWyD9V04o0+60gbf54nQvPBpI5Ge/nwg9mT7mmhv9cBxQfp4vlacnH/tE5k
x5+H0mj3cNBJ9s8Dyifh+xIbVYUi2StyNQyMy2HxMoLW16hBN9KtHs8eyxAezxrp
TYM+lpcVhnLeAFbZer7Qqak7Y3R+AhJ1BsWi+eutE6j62eUUapqxiam4IQkAflxa
i908AIK0DSbxG6+DaXA4QWUG8B0ptTMs6xpke5Yj+T0PUW5xSk/x4SEy8JvxftT+
7/wkvsMhp5xRlRlClc746QqdWDaUCqwniThiHwQUVr39hDMRF+txX6ZTAu3IzPrs
WUTvz10Iwc0uNxO2ex4tQRNAS/Uby04d6uB39LKvgHvAZdFKuKokYfBDGfc5VYG+
/5htTtlJUUu9spEzodH6l+pCjTja0lRsxjON1Kh9e0ThpGw3zlP4g/58yedH+zX5
65HHOFGGL8N5T+C8Vm9bI2hrFXtaIaGXDmUuZERLZcniJcxiiznauqI6AaG7l4G5
QfHZOOJfMaf8nlg12ACds3nfWsER8QgcD3OXEQjlIwncFlv8NzvZ5YatNM1uUlFq
ERaabYp3pnHg57+NL/k5Kp30JlT5NUQDL+PdNG54Uphb0IJ1S19c0IudMbEgy5Zq
G55H4GAiz2KyyE7n+KP7R7omGUlDevQTtbGzEhj+nPm2qz+DUo1vqR1a5zWgkcBG
hEShZzu8pJTiEEHYgXte8hi3wtOMwWS5lJKnPSNiOZIFSscRsUZRAR7vIZdCJu6X
N25Pi8/lxkHWWjHS5L6jeYHoRKSisOoMRXXXTELuGvfMGAKgqehmoW0mBw7JHoHj
U1AXvJraVLG9oAi1Y0C0S+atJ7tSu3+UYj/42HdnHMjmQduNWvj79IlYiBEy5PH2
IHIiVIak+ZXLiEwamMRhXw5vyyJ5f4ppzdQ9Z4GqIeusivsk2IZ+pilxwyw0NYHT
vGAR486+sqKEboZPuYT4RBO5u+jHrAtsmqm8e+w1wI3GhF6oPw9s22R430bPh6fF
X3w2HZoDIoE+2dBm/+D+tZaJuOUTNp0tDBk2MSdKU6F0J4ysV6W3LElwFNkF/KRM
ivinWSa6f5OxPC1LH/tWhEntmlY2UcHWATKsZteeQMEKSwxPEU/lVVnj15Xw3Yjh
kCdsrgpISDbfnQSCtk3LQO80ioVZqNF04sepjbIbwyqPRCMmcOQ3XeYmIzjHR1C8
/PvNPOSrso9Qv5emUDP2EwJeGW4SBCoA18MDA8QIN24ce/gTeDa4/3WGcb6/OwRw
dzO+OAhDeDR6kBpYBKbSUA6MLgdxks+pnaFASkFHCsI22jVXtyz5O527vDsZQAqF
r5dSuuuSFPWDt7Xy5jR5tyr1vNVyYxUvDLx0ebyBGathG6/+3qL7PIisDB4KwFuT
HpTc/udilK8FwOSqcjam8Ze6rx47ENN3MtGkYyBIX1Hn+pyQCYadIFz44Eu4ORYG
DZt9MxcKYbunsRVrDrT3Q8/t28To9eVua5+1CzH2MeV5OWE67f+iUttb7wrpy+Tj
Pb4K34qlOZ/Og0P9DuulaMUosC/w+baYU+Dj637tsVPDEpbJxg0IB/nNyELR/2Pn
oQ6DeSkTroelLyeRhoBjCxb/kUK2upiEGz0cUxABGLgFfVKP4ENEijTt8fKPyhto
4TkM64MZ4jBYlaglsRLLf+9jxXixxB7NHUuFR9FyRKHsowZtx+7ZTbWH0THcaXBw
paWo1GhDO5mARlXWD73KsXKQ2dxQDdvE4led0hLWh3dx7Gm575P6eqBy6YmMT3Bj
gOsL9SX4mozEhcSTB5/S1Re87BkJ8WAR31/eUcbrzVHHW8LLhtX9NJ2r6Djbgnum
WKEOmN27bVUetS7m+zQBvCRPihK0axVjtEa5kuKxMdB/Kl5yNYPsyvN9dct98lbS
SCdBW52F3Tget/AQtpGhesgJMYbe6FKculYBbkWsvw0y2uv/6v2rg9VOv7mtiObR
1R2UNElxUEWIONPtoAUzC67WPwuRVAqvVZK8h6vyVsFQfuVsLEA+mHZCMI8OyQnM
YP5YY3TSqp4tSUlzFL+V2rvce03tQ97kLOy8nhhC9b42s5SoWlpohta0PT8K8293
8DDCkUs1zKmfCjBLFZcfK9KA0pZRqbKTRvtHG/wEHPsmXyKhFZIoqGa3vHb8rIX6
XXnE7yT3BUZ4VbHzO6mXC2cPx088fqgco+DwHOTSdvXUY117a7YnWj3k81n8s9oB
qxQ7xsPVpx+FbV1RRFJfr+vLWhXM+4QySZ8fCIg+ElW8mvcBgs9QHaso8yppSzco
o/BDSCDkZ6E0+1nQq5QvDCFTOYQDgnHwf9sOo6ze3xzYhN10PJBINkBL2syWsDxP
cKnCwEu5Je8Iw8fZmiITDi7B76D3wZHzLBhL6otDp0YVJs+hp77YlHuGwpDUM0TE
werShdhgpKPKPi/UWhxpTw04dCQYdqx/5KYt/Wt7ZG7vjqbIRGvZF3dfRvYa81ci
b0Dlgy0CmZS4wZGROq/r4e4OvoDZx6t7NdJhwzHZLuniV4jweDGCcqbsVjCxoMTR
CO9ivA9HcK09bmp5uKuhTIUldrRfZ53lm+MKe2e2vR5nWRVDSCsBR864Ws9yf5LB
S85447t2cLkUCTJq8FStvOvqUKn1NEPlTdSxuG9E9GECLr5+pvj1VsXjoAjuwClc
k2BYfMiUeBaLB8rkYZhJZ0w6PaULmrbsqW+fBYOEkt7l/6MqbEH7sdPxtiTcHbH3
dlOR12G8nGWGyYHIk5+w3RlL0uKiUW4me7IxXyAP5/7miWGnsp4CSZJmDo5kloCT
m/zGJuKQ+TYWbNnnRs7iWFCu/8zMEZ3FFo86fRe4fIivPZRC9+jKxDvp9gU++IzW
lV59MaYV0lNtUybLe0zAcjBizw1DT0V3vLmkX4K9x6g7+x7op80NKW+otmnfnE7E
e+PUQu3tXm4S1MfdH6FfXK85hY+LaazFrJl7nXo9okhuI93yNMCprba51YEHJRfP
/Ug3pmB6mDPZOOoPaW4whILS8SHQu1fRZQhVCXfacvj8pw3aM922CQPZZer6Q7VR
bvYxf5/PUHYCcV9Hq4EhfEd/fX7xzYxZPmRyAs7ZlFPxkVqliKERviPlC0cSWd6z
4vVYNmixHlBC3VdB8K2CmFEcBuqsY+gAf85O6lD8Bu3SU8wLXilVy6sUw+A7jDi1
pZ1KfxozG5Q3PYuHZXuk60MO6ZKZmdT0Shb1dzVww3jsy0kFCOR/CUWkXCFUfyVk
rgFAlOPclD7PfGOnc8Qog3+Etk59osEnYqH1QS/j42JqcW3ixZKx47LOnpUFVeR6
yKfaa8dVEZxQQACzGBvmf8XLLls0sRYGNCqeRb2CBzri0jCOb4Znz+34z1q91D9d
jgXhB1V1XT8iXaW25Bxo5xt5lZPxEPrLzKoByCWLRWobLpCCclmkCpfR9uq3frxi
wRShUjiuRBPDQcE9igPPQYFED4XjbCQyKkRMiHZAkqzyH0DzCKXP0rlPe0bkfC8I
gk1/K5zBhzhw8GBkpUWoNhgcAHpbeKexbT2RXlw4KZxcxxsBqb5E+9xK4Zhtiuol
XJ5IbDMSMkExNrCnhAcg1Cl3dLviDp1icsSNcIWlwoCFfxJsLtBS4/XBTSCzByyC
WEObGLckrclXbUbFx+hRcgzT8gRmj0CsjUJ01+Qd5S9nHAZPT3T5O+79dFQqqSd6
+0+0g8Hggbw6jC/JTnj919O/xBeFO8XkK3tJ+FPJrnSclUNl8PmM3QG55aeFu73X
WlCHOU6aLw5gr7qBXVQ+fXDoz0zYC1MeVrlE8BECVjVQMAIutGm12h/wv7mlenc1
PTeBi8nhStUjZgOe5rD+TLT6HRKvoQK/0XbDFnEMw+uZ5ebXtxuBPXuJOuF8RUph
GanGBjWb57Sr/lrQmbmwpLUe4aE69jtm6JWN6aULBwLCD9kE9w7VZf//zRUNfytf
Aco2wJnpaZl1l69CihtTmyXdTf7SyKzyw3UI2n/yq+RwVCf4EJ1hKbdbYpRu8sk6
JW80cpPzbuz/n+epqh4bjsdzcmCcBMOPRdCvK+nwXnvbbvTFFwUJILNMWhRrvfOF
q7kU5F9qn6eyD3vXhd/NL5ehGuAxuZgaWGrnzt5cOefPwmCtcR+C9a0lOuypyQpp
kJBNDsgCSTELWGfiV7OiVWWtdsn6wbkWsc4z8PtTZKgBCWKhk5y5OCznnV5kDzqM
bYN5SrvKNZQSLQQbezqsLqhksZd/4rYDDz5Epx3810i6b60//XiqOxevZtLGnlp0
XukIqrfF4r3roBiTJpFbxB/pBwkqiRJlPye+v28VzMh3RV2Qi0Z2NXjJekqcglar
Ml/W74zh4gkhCYQYqXx8tmaAT3QnTo+86LiGvtiChV4/48cW+dNSp1Q6m4jbxfsI
Dwydx5/j93lUhZ3GSl2EYSlQcyWADpFdwk4qnCGGax1jS5iyXLlzYNg5EKbdnvhs
O4Oo06VBn7zYbXDmAVC1H4uPw7U9393uxbXWB3T1CFMrLVFO76YqzLCY4cgo92fu
Q0cxgj0X3pvm7cU5ntQOBetNq+SkV0mLkLWeML/kfoszqhPK3u65+/vNnLiGpqsD
lYo7oc22OBGz7B4y66JN9mYZnPVErHbEVIx27Nx8m2TXWn0ol/j/ghZSeXF14Tza
2kIxTKgARdk6gkFD87Awzdng7ltsFrgwg48GOA3P8GRsRJd/8Tej5Kq7/L991+V0
+8dzTJqqxgG/4iXMJ+R7Hv1oy5BJ3UI4Hwi0Mq2PQIEchRnwMjl9dl/v5v+UXWLa
3NyvIzl0+4dAoC6F9DRKS2GiEQIrWZPUAWbpWtdjEJibSilZdG85zXGYtv8sWKzx
8pZLGGedMkCaBpvVeJum5QP88T4F7H0H3JJj+IO01oyyM35Tnd1q/3GPKVIiGh1V
MmSG1Y+gxrqsYvacPDiz1lOfZj+BBWLPMi1D/KVUVVVG0P93mb4BIau1KCa6uydW
6vFkNIJbaLFxhnsh+F8E8RFGW8NmaOlq+jBMl+BuuJ8Q/4kcXXm3Va8lzApAUCWK
4uBvSxA8/0iCoKMotS7N/Pd8y+wv5PHkroqQSin+QVHtXbtcNCtumEZN5eLL7oIG
y4fm64+SswZqZPY92eprZJ91umAnEdy9YQW1flYzDLe61711mIsWpSIabLM2uMwU
bltHZsF33ygcLM9uckj2tLzM8CTYYm9Fb0WMjO52/Q7BLxfF7po1DuLFLGQ8vrpo
mQyK3IIWDdvj983hoQHdkNSqP/4iO8TXe+Sxf+QQsq3eqpF/so8sl8UBKJkgLaqq
PFSMFK8gTsAI1bYOT3/GpDkrE2rxBaqHebE3+572j9zr3k2Wj5EhrGKi96fLeziN
UOl71l9v9LmBLz5KOEYan5HOoV6MOR2zxKp+w9LF/yVJmub3AkjCb989kh9hSmXB
35Rt9SiaFMH0fzRZDQ47ZR3RDqGoGZaM56Jl+lbwFBzjoVhzyPTPG7CPRZ3Mp9ja
cW2cEY/UJkwhbHd95OV+NXbmVgGDW1TtmGo3rpBGjHMJCNbXrjNlSnpNHebXaS2V
VzOYzmrVju+ueUcZN+kua1n9IXTnIJh/o6YUSVz+oi5u7vKHce8ydIh8Dyp3tP32
7rmPTogr7CNauYQxT+oIwo12qd+2uakIKDnlLnWGyYJgZN4n6ZN0i+TvNsyRT10n
LtaDJm81WkIGeBqc3YUfswGVNHRAAdS512PR1ZlIDJ0dj8TUnnt3QCljdRSXsWwP
Ld0KMX/DObQO1AKWHdlnOaQGBa5Kymb0z5076+bce5GucahjeGxRW4Ze06wF6lvA
6Senzai8iruVUVroFOCkA63WmJ/pewqPMTxWHN21Ar2+BiUd8Fz/e1u56kZf2inx
AKhP/0bPvo0ZKbbUGqhxApgrLKNo1e0ed1JjaH5nu0fJ+3+EqHlEvnQywOiUe8nK
w/aKFIum2y+PNSQR0Nl+30p9x2JI11L7L/OFNKpCKjnDUwxtG3Ezpz5O7EQXUMnn
rC5QLrxckUWOycQ3pATd8FF9oXTyZj4R/xemmRD+7Kr1aRCC30X3Yb1FfkDdBuok
aTsdvlCMAR/iS7s6aF/yIk/2gkuOe2rVX6i2Ayg+zyft2TEwuLDtIF3mZm7xZrzI
8hy1nTdOjm6tLlUksQ99wK+OnSG8Ecd19O4VTfpfLNG5MKRnuV5coAVcQsrL+aPo
LbRlwlnD7uobZv4pM7B9DnIIaiaqcfgNwu/dZw5md9x+l4gvgUpvnnfQ+v5LatdS
uwcAUSlbjceyqinp8V4vOlgJVzNifoO+2WBSIcELp6fE3c+kMLd44M8FVGTvj5YP
GNEhU7Z76teMefgcC7uqXiS233xPuJm0UFYhIORf438If+ZQeurgRQ5Yc2VLsxJ/
tSP/J4e4/s1SJFqGF72/8TNpBWecHzPANo/xLa5UJ2nfld6Xl6gaQN7QMabDaIDS
5GEMaJgkNS6vblbqQYM7DcjNF0ERKU98MbGlVGAdrWDm3tuYeyDaQoM0jAmoJzt6
D62ubb4Nrw7MKCVmpgo8KL/VrIjL+Zr4oE8JO9/2utWAH68Cg//44UVZhFvgefhM
7h1lgEO1XHAwqYZXXUDtC+EN+tOtmPyPSgJCtGSdrzKJ4105YUUAFdNH62Nnqas0
vzhrfIf65EqwSrFmJEQMM9n0fEecVZCm9EYKBhpgigXY4aLpYL82MpBE20CY33j6
bEzsmbw6kLk6zr3IsbnEWB8oUi9yD4xQar9ANEQjI2izM1mxByslnJ4XVh2cksyz
pd4+GodyPKS7EV0rnx/Smjn+ZwvUhia0Ba5k1Xj56rUoN4k4RJJ5UWJVPshHYRpd
wkkfXmmMmQJYY9Ncb2sA7MFoBLh5ej+BCEDlmrkTfXSrQyUHnY/zzEnZNgBJMUi6
PFq/y1xKV+F5IMjXNjx1oR1F0bDABeVal/h+zQfF5pCn4pZhIqfLT8g3JR4uOqpS
3iOxqg+YnGuGs/yxeNEV8DSoN61fXN/gLOf4pB9HV9mXpyPzIIUv22ivqBJ9x6VE
dWe32YPXhYheJDF7qkbqu4Pm3qeQi4jDr2AGJN025jOstDJPQ+ME4sD/bKI2N/N2
iVd/M2mrIC8atmQt5hAZ8AeoyrvxkeA07L4arKAgt60rWeliA/WqiJawxQztLeep
IH+ASYbNhmvHZVZP/Js+A21XHsbzizesCtSg4nENrBIIv/CmGfM8gXPXtNCaYaN1
Ci7S0ork9ybcy3ShSh6qnEowUAyJPBoM2OQuORaPdXbbyWPrmKFtQkH6bXXK7opF
gjzl3VxvaHuZNOZNiQhdRExaGPQXEvlNHWbOlgmkjqV76K2GuB4jZ3LMwbLjexiI
Gqrd8+ylM1G7AyDeHIN8W0D1qYAlif3nThL9TC63Gwbss8X84247aCbBdd/e2DuF
KS1JT42dGMxSU0nqBtxQCYL6l9nAaI8mG7RLd8lZksgOUxfU+qIqOZHCi0YimwlH
RYBn3lp+OoagNiqvEEulZJlfYEtqdjvEupmiXFNlLPa1lr5lnDYTUivwaW3TY92t
uQOJfPWLHhggvfKEZFY4fNIaiuZ3Ne9S6pnKLcLWwwS1MFyHxW9Lksgsu1f/AOv/
jPlqkGpVncngoeFDytQk8aXbC7va60HnRDdO5PsXHljuKJieXnhTwzGLR6ry5pWJ
jme1oQ8xkhPbsELFQ6nJ6vwZM8l3OkP+iy8Rf2WsvDKRn4zsEbl3bjb1sKqHPYN8
YhdLmIXt1kXp98EH97Dby3VX9IvnruLpPt2gJBqXL/h+CHy9vcpidJtd+AZhLshN
c7zRhDuiaDMKeZuBV4XBD7zuGP+k8TZGEAI4WaDExvtJ+mUUUC7Li8+d8KYxlHMU
CjIuZTdIdXbDrQggMrl6/IEbVfPfMREeQmP08V3fmgyS4slrt2sWgJgF2YvgPAss
J+fFatmhoJc94LvCVxvy5VYxL0pcruv0b3fPN2JrXfAG8L1jLbwJVxtF31bM4svf
8EPCFum8HO2A/C5Bs9rrXjcTJ1JPzUoCfPAlvcmgYmglQXZtV+/noyoLac0QQ/1p
pKXWCCclkj8V76WakcU3/uvd3CSKIdl+0aIWKSiYq9/nLXeNIbLJ2y4ZQkhSjckV
6afZBpctfj1fv0V5xUB+y/onfp59dQM47ALrWQY9spVan+nSq1jjLdsVChJ4B+yD
r6HrVKpWCOhrzmp2nKKbzsxPoHCfwQYSaRvhhPPwDaD9JFrjxQZIx3iBjzJbPEd/
YvTAIx2JRNdggNnGefOpUDuXR9epRQlVSxIXzsrY7HlTMOij6F/1F9jZePhmrb02
YSXjx0ydI71txRN862HcLTvVCQfU0aMLFlDsGsu76urMP7A5YS3ALDfn0pz62Ozv
/23mGKiPfIXw0d6fcIOaVLtw4Wkt9O69BJn2AbJSM26LuQmegJRbcQX6UwbAQhbI
zmybvxZYmpJUS6Vg51yVHedrjM1lpW72RJX917kbIAeNj1AhQ2knSJNNuKMOgdF3
+KooqNrvBscSXQUkZLH3JM3twtyPKRWHdXzMqjpKASkuKnvX8fLPpYFFckyz42Zm
uktJ89kBdidZaI92qMr6kvw04c+PX//UJ46maBqOvIy8jSWw6rYz2mbvrq2X5Bt2
c3xJQWAENEoOxHfgUMGVTdvrz3vaSfvIRGGQPV8q6j+HYkMOBhph1s0D4SJEgpOn
5SWV4gA4VELGkO0bnhj6lQwcQ4gsfzRxMSpGrjhXk7GyJxwz791vsule//u2umH5
v7UzrY2wpVZ29v29CRUu9b1lkt/70N1c46y2Q7fy3E7ZqZNSC5WAXn6L0gE/YFRb
DvhlAOIyVl3rBaWOqfBVrDfttDHfGv1iTYjAVjhT3C4k/9OcTzISzKdDw+MKSZG8
mSuc2CFFQjDzEV5PBFa6RPW5OsZG1InIHc/0Xfg4x1Lby2wEkT1Q2igRJq+os4cz
shVSOT0/Yazcn3LtvPAizEC9ki45/Q1USiBB/HSvzV8ekcnw1x+EVqGQFPDmh69r
k27ecuaTu+AZn77So0ElWVi/V09nTUXWQKGBGrGVKhQo1YDEL87gFdtRhdEBf3Uo
BrVTgdQEzKRsZLJ9Yav/Kq4R322WgStY1tWvYm3n5e1Jb9Z++LvpbMiCpHFVfhOH
Pi6/zX5cVM91dPoAvNQE3zLVxhPrJ1114fN0BGwjQlgL9lkyykxjcfX7trHXtMnE
fzJ04Y90kEJ1enmB2fIl2ddE0R7uF0KB2ui5xGF+1Gpv3osp5LY6oX6bk5GeXY3F
ut5sryL3EcZxYQepcfIm5YyYFYbi8OrR2kf/awDlMsKN0e4ET+qoeRTImXnLjEor
eYR45ngsqJbwKxJ9NQixKKqLUblbHAdJzS3WOmUg5sqxVhd/ledmxh9cB1fQvy6C
WFoeRCg4IpXcBpVlbBoT7FN8OR+OmPHH8qHncG13Qbnt2bqQsjulwjnTyftNln44
XIYaPIOr1jJ6ANXL2Sd24VPYLkkTCKT7PS3VHLUYHnr3OxIBy1wpGMr9oz/8omSI
yZhYa6OWFSmZWjGQkbpPX4bxfxr6PJUabrGtdLlw9KjFhJa2T41rM7ul2kq+dyPL
eEl2TQI0vlP677Rurg/B8cDBPvtB3Oh6z0Sjz2h+eJ61XJ6445iAAKUyzPqRiiBr
qxGBp0q9ro+ap1xQUdMeET9WbOfi4+YYOF5NkNit9UaHvuCUfWKK1EC8O0XMH0Ws
lTxbVwtu29u98YbZwe69wgYZ4RtXy325R6HE54vZ/+ukFhKU5Z4U8JePjcvBlnPz
4H4eEh0a3y01Wc9FFlzXRYG13tRoq7/Mpt1j3kQN432TPxWIuTtjviKyTru1d9WC
GqN/1uU2g6aCNDVAdlGvcZr+Cd7cn7yAYUqibiPvtXHq3tMtoLSHuOwNfhl5zYal
ou+MaOkx9KD/ISiwmBY4ZSV+kvhX7iT3kYRv9yOSwOnK8LKXIPNj946uEpKecRUd
G8dwJBPd+bTkkRUqzIhoHjRqw0rpjqPQQPtMPEQsNMNKCt83zzCnKL18cHjDD7jo
SREx51NbZaEGwjWtLN7CDhiOtgPUd0JqIhfg78hNBuv2Oh/IAYBf08LshucQ2gt0
sUbmp2AZ/zJtOKan5abz6sEvShnMdFqQ4c/8l8t/tqsS8yhraCBgujbBWuV0FLlX
CCJcSfsbm9Rt+hTvIO0tDLl7JQzDEGOavNgdpo+2LpedaAMQee8q/RfCqCBOmbpj
VsN3z+lxRIvuA4ooHi57HWvBN6FEjCVAMztSCfn5f8/xq6x4qjdjvgKviuSeo1al
fdB/01esOoS0wgU6p2g1w1jHBAqsw/BxyH5TRA15xBYkdB5jrqDCrIrkKr9/HCMQ
7tgr4Eky3KQrvkHTueKff5/LMY/knPuejml48O/IpCcpUBaBZ7u/8DfkoT3pBLzX
LDomIp+Bro7nbR5DA5xJN27TXGYRuh4yZvU/uyNonXteG5Gbrj0hQCMI+RNbSK4a
GFBGjKjE8pyFgAraYSDOLJDZ8OxFn36uPtIiE3tz2/Te1rQvm3wkdQ4rLcDmjez2
vHcZBdfuI9IgXuVl+rWRAo2z68GQ7EXKt3lHNllN6lsdaon0vFeLrg3ShdOvgTFF
2S6F5Av+obssTGyJNCxbshuU1bfExHN9CLkRp3r/aTF6diA8+xbye1tZsJNefQfy
Y8mfyugVi+x2q4rxT6+W8uFUVkrywKVHwWs4L4+MJ0tjb9KfeGtkbw1xU1LjYtHF
JmOw+NNIOSh+Q8UQd8It1UH7W2fk3bBSMnKPGfFNPIBpDiAdJrh5zDwdIvYqA5js
67sHOLs1gqgLvegpPsePRn22jmrazrMjLAUtI70h1QKntuQ8ChXH2bcNRK/4/ceT
cUQbhA4OI3uwokabM/nxERrDY3uxw81dl6IN+vQC9Rzuy8Pa/QIM7UYGovd1heK+
22n8J6mnZFpzx66FDLSBfEyhOcFFnLXIAZzFkej/+J6Yl9O264yTkcw2qjZahsxO
igubdDMrFXBCSL7/pUkxolmZc/w0lnBxgwdjOivw2PUazSV1oXA1aikzJPN1CR7s
mZtt+DBZVIJR8V3lpjDVtSB494cD/7jdr9U9l8oxP7Wvs8dNRPinKEvIebwWUumn
Pa3ShCRbZIX53tdx2Xuq1FapQOi+scENlBpJQCSZQsWOAimw55Yjbo+DeASs1SJE
kJCuPf4OuVN5iLkf4AmVp5AWcFVjq4a6HbIg6cmnDXzx/STeG7EHYaSt5fK9gxap
FiKlAtf9QKewZyR3LPnSRaczSadEPyF4j33CiEGJYpcSqrltTBOZx4SxmQVWgQmu
oyZFwyTm/0RgE29hvYPKFU9DZbiIdr5NGSgzQrqWLhYFCzpDjUIKkcp4Kmyh05f4
nMHUvin93gotFn1TKnoufxhhFdQ8OxljggM3TDnIMyVmzRt5yucPlkJe4m9J7N9u
ddkosTc4tzH7JhmMGAbNSDEG7ZTB24raG+gV7u3eT2PjI4U+n3FCkfWntIZYNfLA
wJO34vOoKIa0RIg2xQRbVxzVbRH8O+Jo0kAX0aNZz4gGOtUgi6njuLuUszLLZ86K
MzXc55b+Y77UHDFL/AfslAG4lroZbhX/JmRgGnJ5HtuqnEnosf60kS7szFH2+dJz
ca/gxAiJLtboiLJPNJ4c2K4ozP6gFQIAkeIr47XbWMoPz+DS5DSvDdKb4KPZqgVL
jDlj2aXtNpA7mr/BTSNp2vwt+HPBZCDd9ikfbn+497Zo1xKg6cr3qmCylVc3vG1N
wDG6t+zQTvHXEPT2ZQJ1+R/wvNgK9EDuX2gmGE8PbcBVZaua18ZAzNwn9ZmshjBo
QTHHU5K9dD2CM5HEebIeKd5AEmpJ9hsYYa3GUePMiAmYMibEkOjBObaxu16t/ZLV
tEcqMJKgZ/9hhYg36tnq5XbapXNGTuqdchFHbzg7T0lfmq/fwkJim3lyDFivdj/S
fHEo0h0ta965HDz2gQA+zZz5KJKF92AyZMn1NOCxutjCuu5gexKHaqJBTXl6I7Ud
ttpjAZOXcRp7sCQCs4DUjrvnRZ4zIpCtoA96+MeLWLXnQTSCUlhgWCKnjiphrHON
SuhueBGP5ozZe8GfEBBnWrqjqytGJPnXxN7Q574R9EotIJaJwrDyPAILdnHu66jL
97vF7FTeMqFCk7mqfnEx7jfjuCWGw840Z8TvxBnEjboLLv4tFxtEoCEgTkI3hsUS
bVelItaCbBt+kxyZzLC77FX8qa6N0UDNoyaeBxhl/8VeNtMWTNh+uTT+1n8ZC/gr
Fz24N+C1BnT5hqmnIQMyYtWVsz84UzPe9ib9EDMnfDQXRe2h2qj9szuXvM50hzxt
sb9FB0js7LOYd3NpU0ZJuOjp7I13xSwGcBaRlAKxG5zhvJ1ZbKDHUHAz9ZqE3u1v
jzBH6//oJ+piY+2Sbb3N1zKnZ6XFmQ6LMy8JTnU6kVpE/G1yOy9VK9KAEXDcNlzr
FjPxeNr6ro7XhzkbgZicLSC/ct1ZrtRveCTbHzAY3FyBGk3GuXWcwWJ+EjJURbld
s1MhsXRBLfarABkJHzPKeFyjlvYh3mT6Y8RhlvVwa96gs4ARoV0O4OWhJ3jFU0k4
sFhU5xXGJ0ceX/XFh79q13hgZv6aTnaeZV/M8iNQ/6JIVrFjmEEIc+c3X0N2i/W2
CcBd5QT8pfGRJL3fu4arnHsKOOTJ7nEbGKKnqQfHhNiXJdXhmr+qixHiqrD2wn4/
wCyyWtkbFJO77Z9jyTritgc6Gc2dNgEBmLaSaBxDtx/HYZtoUQqPfXl1OcaPJN8z
sAaY4AlRRV5QU7aRLRRnrWKKHoV2OaTmK9geLqikgr743z+/9SLCJUqT9/oMcGsg
BqHVPScEiyyIQUn4VYwUGzFGE6Noll9ElT42Q5fWiGj6MhNbSv4S1aJhZjnCsb3t
Qe8vkZuJaI1AwmtDKe3qfkWZJFqP/U6xU9ZrVWGQVjx0h50PX4mHqThBLmJtqXdF
rKzFEVFuj8iYiVFEsy7+2LaY1mo3yutaNJ/tWpk6GB4RGZmUqflI9ED9z2QH3ktf
0M/c0bPuEjofzY9Z27wMN5R2Lq/xCFYfLW0X0s5irPsvUw58XbTgZaIru6agKkml
UL3OW8FCGH9yqcgGLRCOo9zNM4CcZC3iWQ+FnnEIwXbG9s2G5jJTgvYtwq606H5G
y28h1KuXp5nDuyPk06zm0ZdaZNyx3ItPuI6S6YodLUx7ya+c2sTMhRwZe90aJdti
sDVcG3qo2vxaUyGI1yWRN6dfnCCD35Ub5uyBKY3SLuqUSXVWOxP+01zas0dKW0jB
Hi+kimo/DzQPLRI9a210L1/7GsTp1VlfKVdebDTWBBQyERbai9WFUXahM5OAQrj7
Bxble3XmFpf5wUNd44disBUgX+6hNQEwgD2BFEA8mgJkQdLGAved1UJg6jJ7zllo
hOzl54Pdxz2E502znksnuf5Gbq3stMG99zrh//dKr7L/skZ1x+41FGhR0by/Y/zN
PCzjpN2nQ2TMa6IFWN3kjrIf3d1uPFo2q7MyRVm9oUND7enPqb6T0bxn7v1Wa50t
8BT3xfCNUe4zCW4yzMYuW0mKErX0SST8QOmqaiYMMP3fZ0tBjZQGZh5BQq0SbKu4
YEDMld6O0HSLmBEUUj5pJqgnHfBlbM/6asmQ/n2vXMMVhrpOXrtdLKHX6Eb/ufq2
Wx69R6Ei5UCB+BF/eYPVqqXam+sSO/GPP7FNh8UiBCQs0EvNnS+WTZd0JSbO0AN5
9vSgiwiAel9UkCY6k3EpCCxCnK8z4Wg4iIbNMA8emadmgoBdiYpQpc1EB69Xur2D
taLVSbm05nHWyVLzhS/iGDKz6k9XoPrsakOb6QBooXbSCkXrFza9B0q2dBSSbEt1
NDRej3M0ApYPFvlWXvigoGVM9fvDqc89/UaUTvhRdjdzMZzJDRp7YAOaQWcoGsCz
mO6zJ/HMtVD1rICwWfIdwZc/KTV9A/XaHlvFLYggUDgmtuEjVcI4GyNcT2u+H/i6
Vi/Ym9yTDLrPk9rEVIh7YAkZnFNus5cjQmQwyFhYQERHBAg4WB1CDvSbLLlpTb1W
h8PO02QGz1O+Do2UFnxBAShmWcB+4FWQY9Kec2OMFgDDMjOHB0IWq9ljLuhNctIY
XmN6M17y0gMCXvCbagOGQSxVC5wbxzILN1oJDpJWQ9F5WLb/c7lyUKvDddUFtnnj
+YxtloU8LayqVkOkcPAQimOZ987w0/9vhpM63ujcs0huDX/Mmkh1YEBpQTLnxzyX
sOgU4Jp+RBdc6GEqp0Wh5I+OBbZQM4nGnnp2TtrqS+eb6hxSMJ+8zuKAzkX5ouii
ZCQVV681X1GwJJgzdsHcOad0j/pe0RT79QcTKd5qGVK3mSx/TsYIZMiokDhOoNVr
+VVXI+cNYEwKJT5LZR+efy18BnX7u4evdiRRYultX0s5GHxzCoFSTnPZYNWCY1F0
y6S8c6EseHIhHBObQEKb/+tSxhCHg6to0xxHjK1VrpMSl8w3V87PN96zWomkWW0Z
dpnaBBhFkx5t4wmxnQUYz/mYd9rq5S+mzqRpVsXaduAcIEfp9fdvmwhjFH4GfAzV
eiPv/Y8aUqbsEPR/8MGM78mXbjP+ll937jwUcW4TKEEZFl0Vbt0s5QkR3zxl/A7R
xi0rJVqWEGLHuBvMQNxYiBVsz4M+vw/u9snEK8g449dby7rQM55tLGd703qOEXYf
qwb8IxiDzMiLCd54P+uqBvHVcwUQli9lpjnHO1VqRRtIjhxzxw1bUHmfj5A6gwJd
+K1ZzNuCwojFkP1wE+icIIAo+ccNKQTYObnfUKJfRSpuS3AAPED1sQvuSPNASw8S
U6lSONjufoJEZF9KCmOBusWdAIgT5gwSoO+YWFawP0oU7/DCYFyPxN4XlbyGBq0k
68ZXwRJZ3/sdVdf9kyBUABJgpWV2dgZe7MkM5htBKZx9SQdnjADHPcocwUdZnXTd
VCdpNRmR7Cw3ICUPhGabWEUF03MFsE1ZsKfzCIxuIfuHU7fNd/HPqp3myfPVeyf0
Rbe36JqI9J36oOLZDhC/qvh22LbCj/JQ5kphiraCgByskBLNH5MGJc1yOt3ZrnX7
F7ogThQHkCbBTv3OGAxJtSUa/j09RT9IdITVJcGRSsmul58bfRIB9jyIBeBUHsFw
wZa3rDsYVl9VXoDxEJ8JIgY/De0xUzmNxm1dJAwsiBri2v4SMwAjzbim2S0XnxUL
I0QEEqNsFJi01O22Dn2PbRJh0pa2WEjM96i7Q1SF3dblKbY9+eziBShIPunTWcRl
p4A0wV4q6qehXALMTuWtUWuG+ctXAYlHorkKpRzP/N5nXhhseiQzweoKooeywQuA
ai7RDcPbDjg0wjKIS5aGxUHYU5qYDU5RpTJcqXd/Nyt2yPf9n/QmROcNO/FYdJ1Q
kw6qxChuqklOkhno/I2G5lAr2py7TPn0EjJag2ZJAwCAQ/pLuJPwLOe30aTEFxIA
HBn30qJvbTInDkh1qeWpEZFZPLALLyNYA1UKPKluyVG6atcOCnEJD0lXMcsm3idT
lvZpLp4vFKEiTZeHQl5PMrStUaAVjJbaZTJEAF9HyTh+5k06GHSfMVodtkZh1HBO
NaYSKIGbgRBftEUhLozx2zu6aMgGrcdVyMywkozsuu3ku7ZriQyl5iFFg5pMUOkt
64n1ytcHjU8XBnjR0MX8WMJ5P4bCEVi2mCJT0MPAHOx2YACAHYSAXLNkuPurYJBD
pREs8SeQRswccMmh4kQraIM6qnIkHOroYGzf7wDJSqhXj5Yg2sPJcVN7jnWfzVhY
8uasYZpKFmfekAUTlQu6H+jshAq5Vjr/Nfo1VOprByZa6fBIWPYZg9kFpqO1VbMK
AXSosyNdZCkNde5Ey5+0IX/Kca4RdCNoBuXZ/L0Cy62FQLX4TcVOBhAzrCfVYBM7
Pdxz1jDTe7hC84Dr9leFcrcQOUAt784ehq8BX5Z3IRW1EXmqyRRUUD47JwGAasV2
gr5bMSjJl9Cg4AHtdTYlWJDqMkfkR4+nDGSTTqEKrDs4LUK5mjuAV+07OoGXyKAw
nqDeiUx9TvCxV6mb08CAy/b3TKEhZuPpoY9Ee5XlYc0N+IRyUW4mRj8k1KXS3gdV
009hAG2n6/hpqLWtOJpyk9t53b5X2fkTMXzVmVeI2LSjq2hYbv4UTUyiwvYpnUF1
696XAqEBYeQN6cHWPDcvwCTp6qqCtqslfwYtYcj0j2VYS1HzB0FrhyQsEIFGMscU
6LsKo0cq4W9gBCjA1yDGUP+az4vo+LqhHqxclYvJfW70kMfIvWdBhff2xqiaH03R
YSgkFbotKhew8sKQtpVq6f+5KulqhSm/2O12nghIkpmP5obORUtCxnYTrioDkD3z
2vToASj9yH7JLcG7RyGObFfTQDGAWxefUPf8deJqaNBX3A4QU7K3aUSJ1SN0HqUT
aEGKBviqB3+fZ7ZKrUXKk+uY8tuN/6nvncaSIeqEEoUVsivq1dbiXpj02WxVIau3
++uJovA9+uz6oVRCaYneOA3V/g9/RVNBaE/SFjL2zhQjywF4iP6f/b7KwQcdjGK+
j0FPCCHPOt/JuVErpZd88EgCy8DBmdFNh8lMz/D1JFuu/0R/sNfhQDInQfBy7eGm
+UD+oy3TNOnoy6Q4EGy1urZK65Y4296Gu8mNJbSiOE7ivY2Llg5Nj/bu5dd0AzHV
H3owx0D1bbkOQ+hWS79EQSRCeR9miuSBOAtW6Wy9vRVAkcZDnjkRgGH3ps1EXz+K
tFntWiseqoSHxPrLiyzOdrpNSD2WSaIt4jU4Dol0cA2gc6adKg6zw+DblzYK2Emf
+7ekqPduUCFNwqGYSkbqJUWr+kvvhfOQjlU3p7g5Q4GObpY5AyNEtuCmoOg6q9mC
vUquUQ6S6PGMpIWoTiJQWMFzszfMaBL8Gn469X/2mPaeN1y65xd+LqHnuyRV1BKl
qEEVwe94nXwUrb3Wjt82N1yWY7kGi074bMbuoYW+YT8vYka6blsqlRAIOaabWnmT
6+zMk903GIg8VXkMHfbiVWTZcHkwPNHm/fx79Jf1stB+l3wTLWwiYwxalw5QSo7v
WRa4ug4ATM962SgO0j46uqZL2FO+mbadqyb5F0t1uMCKRQP+0NE8UfgPdon7RppS
8cUthShkvskP0kZASZcskYUlUTPsCyys14ZfbnzqZEyA0ujmRowoWPaqWeuIJk2r
nrBjNog6nHzPQ8O7eVRXK6lhjS2RPiWakOpLJWHCyGwhcigWfiZi+lxUPn0joVmv
avVVNVaCuf1WoSz2x6dwbnZNyLq4EAcA7F7QJ7mO+vUGNtXu619BDJNHhYuffzzr
TNqLCoNHw+qk41bZkqrzVaOOfAmdtSCQLpwtML32vicC1IYj3VpeSbed7tiJC0/m
zbfRunMkP5RV99bYVDytOEshKx1/CDagXdN/e05DvQdj2YW5Wkxsso5iT8h0uyYL
Ql8uLpIIsRndtOBAHK5nzaYSrSH9u0Z9iVz+as4/3wdHDfGtfpD5xPFPgP93rbwb
9RJIs67kUanWhvLfDkgIJ7z9wfVjxx+oroyjunUsgpG7hrvSOUD9gqAk4CMNQIRa
LjChijzhlI7LDIuENyYKHb3mqB28AqGRTJs7m0HvM3VJxjEe8XQbFaB63NJLHCGw
gitfP593Rv1ZXn9HMT1ZCy7SPiwC8F2euz5N/KAL2YBFt0yytXuRV0d+ocyd0fLA
21ENvsuGoHHE2czXYSCklv9QBJx6iI0Pp3elhaCxErfgK3h/0ASX/Orou9P/iDFA
vY78UFhPLls0c+tXrf+ZNoi8tVWIF7L/rVtVSu2fuFIH+/bKoqRtPysQJnVEqQ/j
0k5v6b7Bl0XHK/e5ivNY9Qu7Zq3dFNUiUXhowSXpEWR82WggJS5HRLQ4tj7eL2NI
Jb3ovfCcfz7lxvZh7vkS+THn8VekrpiNJSvyYwoZrg/5tEUBofa8D5UCqDb5KnyL
mAOJiTcUiqX/bU66BISASFShVyrlIKt9RW5qRVO7zI6PLrHEfFs6FYhPE+yQ3CMM
QFspxYqXFZ36z2qpmSOyuTujsir7E+wPj26auFu3rA169+haYg+XyoL/dFP7NQPm
+ykuqKudbUBT7WYsBtoFnQcxq+XPDNPcS8pzt+McaHR2WssV9fS7eZp4NjeS4vYs
yaJtk4l9QdUzYz7H4q2TRFVVjS1QeTVONsN+KwMDYqKQmbUuog/5M+83cE8jOCi9
Ghixb1O9VJ0+OoQt64wXduBOCtSOja7E7GNc77jm8vCPlyydw3mrtCL+AgTdhxel
jSdm7CmlRmZ3ScbhsdN+v5KzGyC2QNmq4GUJCa9O+K6AyWO5piWEOy3/PC6bnkyS
sotzCqerLs8A+jZd7djSSyIaPc0Sgtz7bup+ISOzQkysVSKt85PwNCQnhUzrIN0v
Zioqu2ppzDSxh3KjEm80Ee0qzLfB4riwfrgQ+bTZu9RHCfKYGA8rhoAkJ6jLaBWC
+8rbSqNqSdKb8EflKiziFsf6dYk02rp6gjJA0cgMouDC2y8r+15RvAoXirwP53Oe
t5L/10gdR40kkFrvzQ7RnBnkWkRQwLszR8p3TD7pBT51O4g4mxnhDKcuxTm4IlDW
40JcyFEr3IHVr/QQXKBqbJCFGTad87dVAVz5eI9X1bS+CGRe7j280KFqWqfgDzJb
T+HbjqtmCW6+fBe/NxhYgpz4XACwmEzNL6SKfac3vbBLOW5pD9Zraiq6axHFaGyA
pEXlOTc2pG+U1KlK0FbtCL7CXRkPXPuCC6jOp8oFiw3HUCKgyy+abGQlRnbuznfE
XfhqoGD0LvSjKdEPw4KNf6GpVRsJK6NX2h/2NzJdhfVtswmfVh3lpWjc6mIM3Pxb
D9Whd2apvWB5vF+7XHETkV13x+PkrNiHXIxK8VkwxBWrJyS7iH3w5iKg1ty/uDXZ
MhdZ5C3vfs0yXgonrfB6XBd0AKUYtb0qA8EWyDh7ZgtevzbEQ7KL7j01i+ZZ23OC
XmxTEbl1bXBHchsttRksSOCRrT/QqfF7bLknKIBnBB0+ody5yx6m/IGkLIWn2M+L
DPXuFk7KRHYNO8CBD7TW/ZePgbDuni/E8G5l90HZSrLnx1YRelBF3uwRataOcf2m
TlZms8s6/o1bfqytd8+vIfixePTC0DwJhEKV+G3vEKZTsQVWvp8npAFpAPg9yovQ
L6VeG5hsQJj/4+wDNEDZImDDZ6iELfVDtplOKYyrgCfbnVLzHxIAKH6mIDI15cKU
2Ca2cp/sVudnzHih1wNXTtXarMsCP255LH2Gvem7UXATqzctKpJSRmFNuhf2DVq9
DtAnbY1hZOShzYwVGUmwl/XcEY9rY9+Ak4MUfyZFR2Spnq4wWMqSCKU1rz5s/d1M
InRFOEL+0Ia8XHKvuAv+FnHlFcakXnUZQLWqXd5GyImhcngELvKP70szhKZvQP/E
CPJuRmQ9hVVkuB4GfefLMArr/lOACqYE7grrqKE0l8R2IHs4tlt2nV7EOI6WpmPu
jBBvXiwPx+dQ+dhtUkzpV3NP29WsVD11O0LmjDTmVnzC953nzmLTJbdRtyf0Ncov
1R6ic8V7DxOjF2e26SZtdrzZmGgymQh8WUR50VrIo7zVY0LALtz1fNI2PI1RGzq4
pGnEcoZxPQyVd5p0hGy7ueBddWQhBjI0n+dqiEqeuhow0prURGhUnYx96eBmr7Ug
3aM93Swk+cftrLzRXexsBb9KlDcfQMLwZQDJE7BWn8T4qiAdneLx2DWdYQ7pgMOo
w2R+WCDLczCwnv8Kfe0D3gRufGq9NegBXRj78Y9u0Es57kyo7ANn4Wz7wmWNWGHH
mILmmStJtnKoS2F+ocDoqf+uhz5B+gDSQmVRXcVMdtYbBm5HADSLOWp+ioLaL9FI
m22xYKuqA7Yit769uvZ6I0CMQTPGHmXL1VVbeqdnwCOn2wm4yuKAl4PrHw9afT4c
E+g9pJEgMUB0OVu9LoO0+8WnuZ+8KuSMihi7iuzTSKUo3AomrZ6DtYltJsUlkH6/
O45mHXjFxardtuGP7NxIVfk9eO/03DgoUIjKj85YzM3IuUqeQqpx2ciLT1H+aMsd
N3veM+dya6btLgPeH1+3Xd5Pk/hkVXdBUxytXSlLbSvUAREyUlk1Z10ajgjsOimD
7/FOexaKDsIdXeHkiGQ6DbmlhxlRCrO3Rb32wx78haEq7OLRGMka22JoazNtpiv1
LjrYrE2tfFB9zACCoMikvWRQG4+JGaB9JDniXa7lKPvXWLDrivVN17ovejqDM2u4
Uq8C3bv2CIxVdmgpIKUOHN30nrwiPn5f2Ub/gw1mxjORX6GDOMoOD59JFmlUdR3t
yUjAmNV+2TlmXNE1gvPm1j1+SrP8tM8vH6zcmSlGYEvKi2aiUsMYZMN+SOx9nDdi
phpnTXDrh/ueC+jKh3PY9yLFuADz5+d1VqDCWf+B2zbKg4DeoOgR8jRZZ5FyLa7N
nwhBtSgRpzLZJSNiwPeemvU/odOi0PNtlYSoxMvHYUPFO/Tj87QahK7TWJaj/64E
HVqJJ/x1a8o7hlbAmfQqVjA+/gWc6532IsxGzklZXBLtQrYQBPUjtghF5r2/T9dL
U4rD0fVM++60owQECMsyKUXzCjmAO4EB+uPPsl3xy2CUk7Kta6z48enMPlUjwp+9
/jRShrAWYeBrlILuD/NeqVxF1MbzWrsRUr60vIc6RicZvxp0rucVDSsDmZr/R/lx
IWyU1GTOfC5VG43uEvZU/rBvngARrSoVjBl3ACeJ3kIcenImyIqbdNc3Bvj+vIsM
xNdRwNXGWBh6lvxtQ0cJ2eQQbPN5cKneuZnpKtYxVAj1OSnuAEHvPID/BZVFosec
vLpsrUWUksHDRuVa8EPbeTEVrwO/UQoNleHnQF7KNBZWvRwbI0xViOpp7fPiajz+
QuZYpq9NiTL+64j/DQmc+khEjRgpQU/I5j4bHMqgJeBE+YX8oHipjtSPvAbvbVvO
5I+DEaMxbPXc6Yvi7/xC8L7cBe2ZS7E5/zz+EY8KzfExbvOARbfgAGnp2EsW8OO/
IQPBIpNr6d4ozIp9cNiTmBezROqvm//e8KR9mFf13S4iXxWZXxE7ZXwqetMjRXAo
IX4FYHm0kMhVAk19FhHpkq+ky6OOMWkaDOnFJynq5yHOxUxBpk+Ji0+/F/adO4t2
u6sBE0HeiDp9+6QFlmqZ/RGF0x6/eOc8o4jir7ghhEl66+FbZNZVNJWlL1qp2JbH
/bepsTefSsG85N1eH+GTd+G+Cc8d+omfbK9UMzmcDM7Pj5/7JX9DPLYN8KwCrXSa
dFTZDGMxaFEgwvVrqIr9MIdIdVFrqcYn9SSM6xGu4u6xuddIynb6g07+eAgLMFEy
vD7OWstdiF2mJy7mxXd36kFThl+qpRhrI51SGxODDWz61ABAA7VZS/PYp6b9dOns
d+Yu/K2QsUwfBvl2z84FoVQk/8X/CFb83sd4Jv+mo5hm7V/FoBgcehUUnmv6ZFn5
ShxavCcJGZSRUe6jzz523LaZ65L3NL07DY7nFV7bVw0E4y/RTjfoJINxVBmt3V+V
YLcZ2gir0EBEGuQpaywYzIOOgwBTp+gdvqTLyN7+akgMkY5H7rYRnrtdrhSNZ9GD
4igWLD5mEh+MMwTMJRy6uSYGCc9UcBAObnFttwBmmW5rXIMS3kFZvWAlKxArK8Zo
U9ZSKaV7YpyG6Chi/LLBugTyDg29uwZ/Akk7kUCcDmWA0fZuQXzDO6a4qGZ3VqZh
5p7FGU+dMqL0cOkOaiApJ40B3Qtp/tJcfbEpbbsEwvOtaXCuircUbr7aHo+E2WLJ
W5BsE3ksbKTZAHF6pgoxNlrSa6OJvdxkH+MvaxI2dxW4XejeFoPq2ifMZAs8qIci
vHVgvMYkxvLuFfZfFmCbJKOzTn9d9ohjMdGgETVsq8cVufLNrvdSato8dujrJt61
ij1N3oKO34jhxUUUzto872tAO531GhJrNIdsg9dEF+oJ2kPRd7NXg7bsDGjPnNxQ
2UD3wZlMHraWk3zJYOYy9iKIdTzSiYbaTQVwd5N9tJ5p52D9SgqkL5kr97e//lE3
UmiSkKFxxvDAbVBZQtfGVh1fKiYsTkHSZP7P49v5SGn10Hsu+eWiCRR+AsxVlcFG
L/mBSvNi9qrFgkMzRJeiYO2+cH8w14t+Fwe9CDPlWtYka7smWxMxk3RhhyTacHo/
FJQ/ePt7aM7Cec7Sv5/cm7uJnbeZFGSftfTdTo8/iUoDOO4N/8betp2rMMfYWuwv
95Jop0Det37rnphC01KWGTN0N/ZWTWdhmLggTdCdnEWwdrV79w/jbB8J4uNZBNGj
nZBvSwtmezjc0dSTkgbEPrsWBoW+EVvByn0dnbpzr3tQK+B3pTEIYiv709PFkKQD
hmAseBKZMlUBF+S0mXXJWVIX5a6bj3LCIdGUcgR5/7bSDtYBpdRVK5iJk2bnqvZW
VNo3vieGrQtVEfPjIJ63qr/JgQfGuAC3LTB5+DVTnVB/CcDwJuiZ+QIzG9kAdOov
HPsFtyYZO+hQ2ZSyBpu9rnUX8Dz3xUwnK99eKGkfQS5fUbheeQdJoJeLy87MSWu8
vmu/15ONuGHEPOl6d/p5cmd91PxiKNaR4SUknxooWdVpmw6UZonldI2EgDV0unTP
vk+XafUw0EB+dbEDh2wUDMJ5w3BK+VolNXtbwUmjzxisyrlFZg3LgZZnADGF59oc
wSY0DFXhw3FVVn0KUdVcGwugGkfc+sRF8fVszY+kNQO99aQMq+xNqyR6xTPm2wWU
ntgjWgOBCOBAanDfZGr8PhD+yvUZ8YzCn0kNd/TN9RmjmvQHclYPish6feknJ7P4
FgKx6cjrb6Tm03nNS4/jJCwIAotR377HC+tEoaJHtWNFm+AC3HhpsbYuXXCq20Gu
6n2yleCHwyvc3FT0VuYwJikQd8lcxqpEjTnTQUl18IXENhQuzR/QeiwTRdoQui4y
ySbAtgFa9kf62OsItrnqfoVVepmuC5hGUvmV1VyByRiBzOrlTlvwhGtyq2ImXQpa
xMddrhOKgbrdtht/pT+r9OTwZDOCT//oUnK4BCe/YChRgLbifg2tbzEFIIKVnwDG
e99LHpJrZuutxuZnygqtZSVO4s3WMGRUyuzlqsqQDU5lb/EdPvZ3GaPxk7SwVHgQ
mQ2eo3MhSYeXGLU49BoqM1JW6hiacO8iuAe9MjSKv1wroB5rpieJWkazR2BHX5fX
2MST0E7+0gHuKENNlhbQcDjYImxb3bhD6Dy3X8VTSD92FUmaZzh5ONE6Fyg2+AYL
Dv8CMJy4MO9iLj6llZkERsb9L5iblWjje/0Qdtdw9y8IHzZg/f2IdIcpM6dkzVg/
XT8K+W6OGJdOC29n9Oa+GqwAYdMy8U+IER1reUsqFD2lEGr5049fUyCbJ/MEVixP
o19TLH0UXUSInaEssiqmZntEzcx8JJtPToTS2wLihF0ohYpgb1EohFpxznx1q94I
H8L0KTT+8Yke79zFCZte3TM0E+hi+J0WNhmkX28zrFcy1XWOcJAsHGXRnoqr1Twl
r2v5aT935gtNf3FLnVgxQf3tFD330V/PcKNLApXjX08DlfR0JEcvy5qYydhFa/Rh
LGXSkRrwopJAI83K/13tG+hUHRO75mE4nNO7+obQOhqWjimFkAyzngJKiEWwVKw/
4WMGY9tM0+pa63o4SLlXPkB5Auj7ysNui7UiI6rQz8anrLFHKVT14qnr7A+4zaCu
xR52N2pul0o7hZEAL0FjtckvEfkLyGI0dkwV8yELP8o5j4GGG3SMspLs5ihWhUGJ
ToJtrR8R6fQePxSiXZdz++8kKOsLx7/zPsDDW3l0HIg+a5LeY/yEErNT8pw0SSHS
4wiZqH79DNbVmJf5dvuir3PORuOfG8sbSB22ppUuffetw0gOPWHdS3n8RPFt3iCa
NiCxoqCAMbcdShfsoce/KhsP7fcaSMY+FJ6/xfKg6DQZM0XE0baUEtcbhr6l79nk
HC/PDvSOVJ6eZf6obsKG456OqSQbutn7H9B1s2Nhd3Zo3LPWPkT/pbp3lRgXllLU
o0yDkJ1ta+ANv+Vl+C5qsf9OoawlAst2ZjsiHwxzlZB7jrGke73x2fitG/f68BL6
/SxCfrIBmVoisNU8x3BFu3vrol4hjXyPbEAWq77TAVLK8TcBYgiNK1bcGsE0LH52
DwArRzH0dcho2AEqSxwFttn/L48ev859FzrJ4IxdJVnx40E+ab1VYka2BNR116k6
oJ71gJl56HmmqhmYFgdExgBIoRDvYB1QfFSuDZFUi0O96oN3kgAGJWyLK0Os3t+6
WRXUJ8la1Jk/F8R30a8tYnWu+7Aeo6m42PPsgMfUhWcnuTG+nroww3wdhrzVz4Qu
57LMvCpL6Ph8ZhwymowJuwczoiK874GqqtkwncycdesKnu1jsCSnx+3jQ7qZeMTU
Fz+O/L/KFP3g7/MiBq3Vrw0gw1Pa9JC0jLBftHH8R9RUSpSb1DfZ0lAaFpjiDGtz
znTE9uGhXcyDOMZOVIBx5l1j+Bj5vmSEN68Pv3qAE0E3/1XLh5IHJhzblHLsRJVB
m/oubmKln371w0b5D/XlZi2uTGP6tY+nAXvDXowWjHjlq4QXkNlq9jaGLPXFxoyw
E8fpvpN/E4kvhw5/FqdiLfU8wDYMXWbEw0yax3vMfwCkHgu6QCGYiR2PPaaJFnHh
UpC4GcgjS4LEwuBchuU3FG2OYWcR/2izaCvRXenrVNzqDuVc0bSusTNgRA/w3BlB
zX9l/9QlJDp1nCAGWbwIXPWkd2X6nUnSiX4vtV9zx4Cyi23xNAmkVTIBJcvHAydB
M+xNS9+6NMc7k1jue6wr9Qx+gv1A6GULSGb8ag14dAeEurKTY0Fc4UiKoysBfgo9
w3bjK3E9DugOY5hT0okdFdg6d+HjCv1Rr0vxNLths0064gg9kwoHIfrF1moqKU0J
8fooNwjeAHXdszFiBrIP9AH/i7GdGyj6iOEIavAQR2dRsDELSFIyuVaWenvrFKoi
CLh+SnxwLhYje+MBuJjBK7NgzrE6EMuUQkLGOlCsKK8SkPs5hpYkzjVVZMDOLcYS
Ik+ZhgIxLIHBSJbzHkXMMH6MuRL8fpgIh+UCH9u7mjPOEeLVpkzCoJgOYWYphHDy
jyXJNCJxbh+5K6OML+etSlmJs8ehKV5DoPbekPjj2ela6gjBJpmqM9PH9VRhvIEF
HBKot6P/uAJtznY4IMNZCfK+/2JnUSSwYzc3WqJmoBA1wu8tK9y2O2QFajAtTm4y
iSwcOUVdJjzuHnUzGi4BO1b6PBJIulTKSm4H25Tmf2J6SHPFffIXOkgqrcJaKExD
SbHwdkKOIWq7/1P3LJ7FR/Hgqlo9vv1fhSCfRJgKsDK9OLzWw2bxERPpIuH0QgJw
hhFky51o7KBCbt2eMVuL+B1mbEz5t1zhs8x3Xjs4rnr9lZsGWtsuUzj5LAyIfHop
fue+oNs4tR1ng+aUyj1NDwNZUAN/BiO0htmge7lXjI8EddBzL20/mWqrLx9H/NTQ
UnpJyCoiAoY942JF6nD9IN5M5lX+wSlYCRDnuKaXFsIarExjr5kfg5yc2SeFOk9W
lXwOTDiM55t1dtUuW88lH6mD1h4asc7+n+qG5YolNDkTtI9mDGEL5LiVC0NfcDgc
XtHvuBfphuQArbt3s5fsg6ho+yjwsfhEp4E7mlkQRW2h37d2isAefWxsdriyT94x
U4DaIWyOTK1zFUpmYlimPS0fNLD5zl3Q+tR+TdgoX9h9RO9ZakwNQELPqdhwtFcj
4Fik2vDAAZDiYQPxk810t5q4mon2CHjdkHjSE2375HZaemfAdKhcyjpQq15jOcZe
al9L9VrdMmP3CM0KL0ulBsVFReKRnSZ9ljGgFs8re03Zq44VdfRT1WTtg2zL+V70
OP6dF9s4vFzFuqiLyZKONZmIKEeGiwsd+93UEhq9B8ZDfWPhU/Wrjm5Tbo3rKSBA
U4E+1K3F/mJPBbUZuqDfbAUqaKkF7QOUtsmoLfySm5ieeH0f9tZCa2gBiADjYObL
d60xpcR0eR8anBKZ3kqJX/F/JjV8CCj2ZbHI9Qax/sIebdb6rvqyA5lKHCYlM7DG
tQpfCkS0xl/UwTnhpXrHuKTwx5RWMBOOQhKlVpKp7Fx+KFdU5V9I8RT4dmeWlJ0g
ZSRaWWQS45mL2FSeFLSaiQ+drYW8YJ8kmJ2GjUBwjutajv8CO3W33gmpxauEQq3t
fGkk5bu2bpwNPk1UJkrJ2XQ3CL90ORv+73HvnEMvyXgZjGDlRmpp1541jdPhnj7J
3nJldhAU3Mnkqy6EcEl/EAI1TIfLY7dq43EQKuHZ0xVJIXuBQCyLocsdsmuVHMhW
cR0kXqoelJudps5KSFSFfa3Ak8Q4nGLj0NTQT0Cj+1k6LaLhTh9EsZLklWYAKQqW
dXx89SZyIPp3DX2OwEHvY2uBUrr7IwujoeJOUXM1U/SFS75dddymMx1w3tJQkkSt
ZoqPpWsDQij5ECB+XpjxtIWKGJItbnFGZ0G2BmhP5ztfVAPXxU06Lt4HZ4rAeWPV
mDmRyyBSDAsSJSKcE5Jwq2l+BEoJHOvWBNsw7sAii/lJnc7Mnf43Wq/fDQDg8WnL
HL/SksUATL992XhUdkJcqrsvRVPwVnPUUnhnXjomzEOvu6s//HNL7lt0A1AhZeC3
Sen8wdHE+/MldWtq3KcHUl7hXnB741KfS6mzmNFZJzwBvMv8TyP/OBirPtiZeOiQ
r7GrGwn7Bu1rSTjhwzbjkwx6paW6wDtjaW00cbEgPBTAtmT6PuhzpwUNGrBP95w9
494sCfo3NqzYbpLhGO6zacWEc0v/CKlZXCiFEhj4nHZXqi5m0oJnF68zxS+6mD/H
wGFOZFhTNC2IQPZIxHJdoLwGwQzIU/MyNd4PcOGXQiN7WtmqQXp4pre0R9zDtHGZ
lRD4Dgp1xDxyHpGJqjPVc/71AJOR4w6xBGGOhekehkpKvd1e/CZuQiuIeCNK3h8G
r8UzptrLscGv/1iXyMizRiYgLt4N6sAB/yHzfYoPx8Vq+31ZgtDkHV3qlOLQpJzX
YaPsun9AD12ysk2AV7xS0f3DPDFzRyoS76V49ZvYhlloWPw54EM07EE9zbmVUsHQ
LaQr0jb+kopckQRtflHky1EB2BoeJcbEHM+rfPBVe+EtqcES/Neu8SHPadVJ7xov
VXDaJg04BaPJqC/0UO2wsKYxRtp6gr10ghO75nCZSoGhuWrP5uD3OXUQybuoMhK9
FbskzMJ1WP01tTe0EUQgTf3Wk5AwT+IlpxVAIaOUideTT1aK3gUp4vfWI8rHESSB
TkN5Wdkj0z+2GbLlUv8pCIImdxe1mXJFBJIOoSZRCWzldGFOOT3zwO3iA4Jy75iF
iXNLNbGD0IJZsHBceVJOMFESr/3Wykrd1IcSnUaR2AFHoR91YVV0lFbkdAtyJWUz
vQ9yq7dMPzoginSnP/oJu0sJjoPOkBINTVI9xetKaOI2e2MxD6wAKeNL1LqrBycU
auen0cuGn1ReqW+bZHkLTd2DRi4qLV2chLaayGk4x+Vgxpt3uBnshvRFZh4JWGf0
0+9c1kbC7HWWI8WTSan7rSfrWXq2h+ixHQjTKdtJa45VEHG7u5arObyaGieRZEsd
usMmhNct5d2s26Rz3yPBLLlAzfwJHYPQuXOFHW/AlUMvdj7PeXxUu02BS/1KCmKA
sh+//cbRIn7+nIrWvbodjJjiHPgMqUYbs4QLQIKKsfHjeMAWlgrRLYxQOiDffwtc
MpUvSxh9GjZ2vX9GQ2s2IYn8H0JipClTm2KQzyH6PQgadkvh1ZPuUM1iUnqbVXOk
jVxxvoAKgfMAesT9qGZHeOaR218Dx9ASRHtRnMJFBmpDBL5tPHaset4TwPBuQaYk
F4VUzBXc23N0nrxEuBZJpS4tJsF098yPu+6KkGlP3XXhkH5fS9sHxfkn98Xp4KmT
9W/6ViIIJrArrLRp7OTsoMVwH8XIoHccoKv9UzeTmYiPGkaStuusWwY5/pkqaQ4p
UTr3K1huU22zCEX0htIdAjRshCXk2kgKzzAtX/fj1G2FR+zRv+4WI709JH+5f4c2
mLRua2i/Y6WpFszrbZA7M7bgWurc75r+SZpvn6EFetm2zkEkfJr7L7piudMSUct7
7yFFZTMSxmYIj9RwJtYIUOcFQMhoyzTDIwLd2sYAAYa8SHdLryeW4V2PeLiC0Riu
gaLALMYL98R6mU6kKxZDZXf3WoqwSs3NMaYgmMtG7nL1c71kChdq5qB2pD02OjoW
m7kUwoFnQ1OoyMTc1ixguFE6Pb2lDyznx7dKTawNPPefZJEDo8G719guYewIKSYq
VKOXsf1asJTjPQUCawpF0OrLVKVqwssS4b7lfXphU54BbIl5gZiD8+Mw9NulaxCH
yMJvdTvcvRiCWoh6KnD7iLFk2WfCERaz+yO2K5UsqHrDih3b0QQUDHzhfV7SkUst
5QV3HBzQolP5885SKhoXARxtgpgmtwXKhdqunwm9FhusCklVVi002lVhpGczjtvO
1zuFWfyFLtQX2cLcxiBQVFccmiJtfSoaKK4VF71H8W8sKzYImn4KNjbYiInY7aJR
bUXCTjC+3gfsa4LOjB9A5ml6hsMQnven0lmrxilq5ze+hgHnM+ZnuZB/rfatKsvg
fVABTfHGtMegYa8kEgU2cHcmtzcdj5BaO6BBIDemFtfGmiSw6orIemQi1qiHIXIR
vhBSqqcNbheic7v07RzOr4k+5NOYjdZklmENqd/0x7fTUySZTIOc/3FaSvgLqnBu
uz+UJEUUbdK48JwlsSRJ5Mup0ZkKAqUYltLNzOsVJjzP8mM40J5wOnge7ma0sWEK
DJiLmmbVblMG3kR4GLwfGLzqvxHaVvg3cyRtXhc/Pui4SbdiN2EgUBqHQVY/Os0N
H/t5RMjmuonVeMPdhAPTjuoAgs1ykVZvxl/VdbPA5LCOOIVm2pFFFE2JI858pbP5
ORtWzM5nup98ZpICAJelfRlV60f77eqAoshkhN90msNugfR2BRGCUDZPMME8IqaI
k0W0YUtd/gVi9YtLvLoURpW8devoXog+W5cIeg7HDDrm5CqloJq1Lu0bM61WjePf
mtZjbfonaEBsS5Eu1WaN4UASzzQcAPVeJF6P7E9LszDI5oO1VLX/W09cFp2huB7o
/whjpVVlxdJWjqYrAhmn0AR76GD19ZBirzFE3zjqfiPr39XJ45r5FfX4gn34r501
pvtb9PZrsfa6+HBL+Zi6D3q/JkVVrjQu4V7oF6HmkriLx/LB8bqtIJFY5VdvvSzJ
R2q/VMXWow+flYDjNOX4Z7HGml3eU7TRCu5qMad/KB8IxJkxemL8D/Pa1ur3Ml2N
qsP9NBXwdEO0jWDgJDg6MuCgrY4NMslQhPvAne2NiAUQ7f93V7s4+GaRjRe6ym2E
RRYtO4CPupX8NXufdmNib0GdRhpnQbCXJvw4poXkpxihNYjEzQ8jkoU38ZUK5VV/
rDe8XTLjvAf8B/8Sv/kD5R/dZu4VMVZM9/6kvXpUjrBvp866oeQWzKXvPvx7A92l
E2k7Eda9k/HgebV1FMkGv+k6PNXWnJO63H6aW9DYM/Uc8G0nrGr3q3mNX6ou24cY
0q+w0aE5W0tNpXVmhzrUtZZfgRkA6nAnZrcqMS8iouzw6dKAjlPYrze+ARssDcpR
FWiMUIgortrfQHllPYpKTn2bgS1evfF1BAi4BjVh7o58gElDFP3RcTRfPoS0WsSl
XySyK4LgOJM6USstzzOupc8U60jy6I05uDZ90JNprAc0k2vH8KW1fXNdc0xnFn6P
IFGC/Gv9X7a820nBUG0maazMdJ/YwjJ3qVIM4XIGC0trgj1La9FcpwcdeykTxZed
R2dBUONpfY/c41MUIytqxHSMoG5lrPKnQ1wd0WDjXzUEk2VsJ+gHRfcO/1rteRHX
KNOhsqfxXorgTVnXPto1Eaf8e4+FFQTiwI9RFs8+p0O0s9fUuA/UncCkrjvXwjPk
0N97GuC3H03hluX1weKRfCW2gZ/K4+1qevPf26yX8JCMxJuUQyvXijxlL494/Kde
Xqa+sXwQg+vZJzQW075ja3+DMGDQWq/peGOSCUCBmpcXIXc/9CADvlXCUTMRUaHs
1hswQh0luC+pdsFuUS2KjL2quxNuWguV8UmcAzt3o6f4YWeDDHIOP3gctp/F/8C9
lLnMbdQN9EOOLrJDcCIVyrPiXxwvKhqIq0PMBi7UWbF95JykCcBG4cJqNCNu+qKn
07h+nPRnm4gLAJRz7txGn2jxStI4WMKxpveTF1Sdg57l8UoNHu4POwAv9XqQe5VM
w9zFQOVTn+Orc55rvNcgeoKpLNQRMnLg7U+XaLpc7lWrYOsxUD/BNOucdeUJeIN9
bxxoov29O7LYa3rqQOAgtGu/GBENn7jdxp7fFqYMnqx8T+okTkjAx+Lv3X5IjxrO
gzzAD5/ystwjbnOxA4pFOvEtWS2OaG+n5eB24IzimATNtwu6sH56jL8Zs8Rruvw3
bTdatepyt9+rf/mNEsXN1ODoNPVK3LRMRofnjqYdubHRw4bBXMBITDWIDkbB96IE
jwl3vZYgvWJSWuThzrYN5G9ZQJBGTDbFXfIMY6zlxDyql8h4wzaUypxLKU/Nr8TM
LSEj/0oN4m3PQjwvBHba3YH/ep1Rbar/wgYCp740LGN/8jXe9X+At3RHeYM4Ra6X
DcVsNc84kRpysY5t89btIJ7IuwHDVVXTGwfgaFjUT/8JfFQEfvr0wf+AuHV8JJ68
4Fkg1jW71ixxzkGS3DitrpPsHg1c6syjwGWLMTvLRncxivTyQ/vK4UiPTLQ+9Tp4
4NGwQfxppey/dG97EoxJEwKTvhPQbF4ydgzCseWL4MKKuMnL3NvfnFtZBtD9ey/i
RKtDLv7o9cqia3Z7mHHopmfTr2q3j00+/eJPJNYcDLykdofeZCfFpBF5DyNX3ngn
BbYCR05kDc+jv1O3FF74vvuw7HRpfCbhqQdOcVdriJEG/tzbQKbjWB7tRYDqfYrH
yxTUaWf/8ze00G9ajMEZ8tfzrvGlO9JN4DJXfPPYEb5WGluz5iHHr78sGAIYT+BV
CFn+d97MxJ+OxTHrWcsZjTfIRxIFidh4qxDbjuSx2RqGYeK9DyGV54HNxCBi0hkR
nsoYpMCnsndo2tbMzI6KpDO79Nk2KKev2+PnTSAZX0IGEvkGO5DAhuCDRakhED9+
ghjjohaRpNMgc9D4b9Asqk9pUalDs56azex6YOhctq+qJfLzKAatcDnZrNeZXLnH
gPAur4xRSQA9aoXGqGve1Fir6I6O6UFyY5fq9dLv8tKsRc22qiQX4DYD5Xi3VNRm
G6umqK0nPC1GPE+Ce2XzCUYreKB0HZj0ezuAzKtZVIK3H7zB5wAcouQw0w1kNRaA
jlbGkqzohvs0oSAbZDIVSXE8iTM8fmJvkpDKqQVYynpl7CEnj0J7Ibp0PT5M+bQy
S9P1DHfO71i7Mxm1sxFgc2xopj+5RYBgCKqZuahfOp+0jvaq4GnfAkETOyrTNysJ
WTBZ/jtSkNZPGnpXGyY85f3SplIbc8XH0of63qzWI5RJvaEgg5hXCBL+/AqVIZwD
QK8rE6X0R4ygsNSmEIzNUeESe6DiP4j2jQS82X/rTacGhqyCPnk+3gmcsX/agujy
QaoJmanv6mFyKbG0alkdO6wnv9MxeSp2Dw0wevS7e4H2LjGyO5POcF5cpdj9nFfn
gKf2NlnNkFbsXStJtgVvhvvuHhy/h5a1O8KyaLet6bkLnDraPtWExpWnNFNReLJF
PBAnktY9SL0FqktYOCZwGglBd0cHsQ02sr8lsMbGGCC4v5uxlc5WcWLKifa53SjO
7pPErLtrinMqlwhlV5TPdce1MrnHa8ieDUhxKud32r4Qu/7PgzSPKZZ2f1kH9lHI
0yGPtCCeBYg0dzHEztLgjIZG3jgBXE7sY15NCi42FiytA/5Os9LOT+CXw5S7pCpk
SwsB7Cqo+ezl2VIdqugprPdojAvVJ+xoyOhbMEBPaCpyWf3wX7EdaM+R3TEwrzlO
DbgHIpT2hVLzxC0mWrwW7qrdAWKGT4I/57RoToe/WHVdlMM9g/Y0oDiB2NIS6CtN
PDVMrsQa7liYLXghG0MsWJdg6ry8KXpOR0rJv/Ro278yrHkx9Q9+5MtEaMYpDyhC
VvPc3F0v5fpIuvzdk1NSc8AyyhFmqNDFgNSZKQfT2WZbPmMy5hrKQ2Y7YICFdFRi
TX2uJLbgaDN7lb5S4NILMZNHheiZe30yy4tsa/Jh+2QmCzKo4cno9uYjZ620Lksf
9T/pGvxb2vScUfp08yK6OiY+YYKAQhscFjP1otR4aCXZRlLrRSKdVgjcwji+QWML
jU97KRp58i2oW+JkRVogMaAIjR6teLjeILnpt5mjH8yh/LpQa4vJncd3N3ITECBU
yTdz3AYpyWSWgXxZDfm5ehsPfObR2uP6U0CO2kpEME+fiav3nr6gvqy/1wSUL6ck
gjROHaNKap2cgfDZ2f0l6+fLirCI0NR8/SKm7+0UdMXggEDcdcsgL2YjqBBDUuGT
H2uN5zIbt6Bc3SbR+Yx7yAwWmt5jyj8Wl3BSeJlt11QouvGULSZpYhn0C/eDwWi6
I0wiYWJPLq2jcq2oiRodcvhiiUDm/5FUBW+RH/MxGvUhjkTzW6YgVo1SXdL+9+fo
R+UVcJrmwYN6IHCk8arkHB1N99VbBSsSf+7DNL0R6wTvfXIfNGlS+2SHD6FmvxrH
AZPLTQaqdz2xl4fvulgEmFGRfCt7UnRYVWUWUxm60GqPgTiwQ4K/Br691PyolgTv
xraapBUWh9Ch0U+4iGc7ITLWL67rgrSFB+Q3vHcCB+Ue7sdFPVnapJ4nV4HEkefS
siB0CRLwGaWTyaZwK6mKEbC2dWdjtXmhncQRaXnW6lmQ5Zflz5WTrGHJvMs9+/Od
uTxVMJheCKPBMvKIeoHgkAzKZmcV1+lhYyzhk6k2s0zipwt3jCOyjTXhopQ1kly5
HzV0Lb6yIXu0ThOlQeMXMGvRawWz0oYPXz/1sHDnwa6sZhf9Lt3fFREegPrKgLTB
nDc32CO4x1ZeiYzzvrVp4Q9dpCB6iuici3ACcTg/DJqv4VPtmcqMCw1BBRNET1VJ
n1Ypk07kjHMgYKaKCrSQ9gBDHxYGuwGL1vJAcpn+JAhddYbmAhImAsQ069/AYNY1
np/06ahHEGAUgAtTA5wamBXxI7vxMruq7iHUAMGfuhZmp86s8iBWxvTcZ4PjBPSK
GBbbz5qBuLal6wmaNd4QeHCr+6gffXiOS/Eg6qGbzf24nw4rB2z/kzVOVtswAJlF
fDnQw5t33r05qqFtUn+3FZdcBgdX5FUZdyvYn+qYiJRP8JFpDrakLsvyOE6wpAAy
U90uBX8c9guXhq3CDnS280ubJfQMafeT20ziSjCT3MP5GYdOD/fkd2aLhkMHo+f/
zgg/EwPZsOyy5xq6bGJUyXS0g3PQo2UJ+G0LNQxFAAF2A2dXXCPsmzjPUsOrMR2A
atRQFUWdCo2oElM7VzTHNf5k8RQwdL4VmQlUtN2QB35i/9S8OvRks3eFTVMp/pkU
6+be6glevzqsWaNZ9Q0IoTmQDha+lq/SIgJnyeygEEwwvTpNO2rwiX/KSR7G/gLf
ONt7mbjhqugPkeZo7eqlVPcGCEGHn6c112+KpJjcVdBibL/aBqdhuhBAu1ka5ykx
Bet/0xvj0DCjcew+thJcXfWzRxJRqtCJDz3tyv0pUzhaMvNb48wuVkPsOFrRZImK
zhooZ9dgZaSaRy2n/A6ilJ7Fm36cUI//jBAgAipTl5VZFoVYdIxqZBjnhqn3tsfy
DpM8QwqddM6tadH3AwIyyA63T1kFbiX1beb8wXOf81ikyylRTZxvFDSizkFQDAdO
ShSnXeSaHqQR8aI9ecppQ3euhukuChDbM6kNdKcAHuuTt8evMYewVLitoF9xdo9V
wIaRYeOoHZKCa/7GO5wZOQ89OtwvdyG6THXoOW3HD9ARp/NwulXqtgM5GUdtPjl8
fPSWvJSAgG6zAqnKrI5PQty6NVJJ9fU8aqIFFz5IKR79Z9zuPMb6XsBZ+0jh7RS0
84UZVOom+3Jxf3wkW75hzKqIYx+VtLo7C8B9Y9O11WQ6bamE5mMnw0NUE2HXkeLr
aFIUSyCQPb1kGgGrkd2NGG27vUGialt8ZL+CjutBfEhYKxCkLc3P0e1atvJJM5ZM
ucYXbSoSOfBplKMnpBgq03Z+LL/lJwV6FsfnVxVgQe+6V7egChFAJmlCegMNEsp2
NoHLW68Fi8jiQOqlbW6qUkFKlxGXyrvmFRTyxIqQWwCySBgEH4V3lQm79VY6AcBw
k6X+tLwyijTr57gCQs/yD5/6fiwfbGl8vWompZLWov2GVVpvQA7UTeq/cGNJrd/q
PQ/sG7okt+LUUAvqQ7U35iIi3WlexL6P/VLqd/6e0Gk7jCLNXmZJOXG6pS9fhSX1
JH69/1YsMM94s6M+UEOnLoe2bb8e9xHFCKSkFrPmLe9jfWCld8Bzm5/+vnHUMw2g
pdGcZM5escgkMN3jd7kwei439tx2jjgZxGfHZg7figfSFjvfh23hD8C2J3C39kwu
B7JPH+XnY1BQZftVP7wdfhM2GJNGEYybqni88VrHEzITaqH9GxcCIvNBVMt/8hg1
FfdI89prptaMPwT/2iVWHUUCdBJul9MyMkMFPWBABNtuHoG3PziYrWoKsJDp8u3m
uXf8yT6bySapioMlIGoQxVbtXq702wqQZGmOSnHf6hjvysANs/8NvBzINGM1IL4z
klBvWjNN1kLqD3xgbDk4AqBEJTBxgB+FlmMyzDMNs5Uy1RmYvwCMUIhSBj04hX+Y
FjKDLqJLn3dSTLDnQFlH9EiHP3zfnf+/7nvWge3S4GuUSG22uBwWTNdnqBmx154w
6ieZrPMxRZh4AXhEKOsEFEY3tDGg7oPdGtZgm1VBdZUxnQxIvOG7Wxzqfh0lQIQa
RhgMAWFmSf5wiV/ZTCASXF2FN8k0tTCmkzhISFxE2YL7ko8JbNT0Nimh24YYnr0G
S1tlDBD32JGyTtdLTWJaq3wmUWqhEMrUQrRGfA0l5PnMT3RDPer718OWrfYNjupV
c4SSF5aAyUIyib838RWN4TTcszg1c26scz5UZmgY/2z7ubC/mvNG/Cztrs35gI+H
VwxUqP8CLYfbLnCH8fvcvjSrG6wnHOTOG7GT4+Uuse7x8Iiyi9zhjApWEUQbQHPh
r3J+ghEmwWbP7egjrqSi7Cj4uSptiYysLF5bJoLG5Owr8AQlVyLm6nazee1ZSAIY
B7KbIIBOfSYVmYUmbuToEalTmawV0+H871TTd/6dytpszFQHKs3hZcY1cBo7fe7y
AEifCzGmyEo9Rk9ZZ4um6sVmM8WlocnTs0x2TnrVZ9IUJrytjjXebhfWE489kqJ4
25wbNM2PyzXOOc8b85aFOCwl5viEbIEnLo2b22w+pE9OEvmdvKm+RlXHdjTxBdK1
i4vWZden5zzgCK1VFGTDLAuraQB/MD8CDSjAiOb8A3Tf8qmbDryUmbxX7nh+QV7D
llZbw2hjhdpt1uGj473qVuwcBJIWqccJBPsdKN6lqioPDAw4wZ5fQaHFdF1U0ArQ
btxdS/QNr6HfXpcQLaFfXzP6AHeBqQrUOHfK7fsYwaMVRAlanY+Odr/n/fQ0aqIr
eCJSOWNWDAGuBnAq5y8asRmJZfQGHzJtzE9luBAI8UIJ4XwYtECY0z2pTc3mAr0z
VZZj+bbPxjU9nMrPx9A2tP+hg5RCzXnprqnHltqjEYWDFB81I7cZ7OS6uQF8kdSh
EbEgDo0ZSgviCkz9pb9xch/H4Zv0lLdpgZc7AZaPVM+JFWZpbssL+RXntZaTE3uw
8ggomtL3eizshoChuvKikdagrZqv5t5FP8+hZ9mLSuc3J/Jy7B540VfkFdgQOB79
LiPTx3Ivg2OIUxGEkPxaNLJJZ08Jz+FAi2WOlcmXI7ECt96MJ3nSDBEjl5eDEd0z
8RKsSWXth+q0P9eZ9X4kRf/lcjRhj4Z091CYuoeQGE3jfETogT5wCeT8rdfe/IUm
yRHMMsY49I5bNN2wJz/vgy9FZJKxllINO0/lqe1GL7IeK/mS28UfIPdMWIuIntRk
SuDBX3vYt7oxjiI2AyFlpufVBwdQKPKn1cpNECxmHbkaIu1JrCGTJRYvBxqlHjUU
NrtT3ts4tvyhKcUj0yfUiMvLXhZWIUId7ewPzIcCavgeI2fZHPgi1UTFZtjYIzb9
mKNbOEoB/eixPdaIcnWIh2vUIJ+ZyCFRTnwivSrJEo0nMrdjAJAsa15uZXVIUthO
85DaebOW5Q9G8NqydN07qsOr4j4vaKStwbIrPooC3hpXCJ7tatUtBcSVsNoqEN3l
mBm+hTyRWFvfTe9R9b+Nlp/IPPoedWOBRmL8PndjTpFWV14+FLV8r8XmywV2SmO4
C80QhGs4s++IM7FXhSssCO0FOitu5T7focp5X3dF4iIPlH+Ynp+FUyUe2mxGTSAj
higCEH2ovTxjrGpIOAVbCfyNfTNFhDAgzoNY1XePxGXzU+6Qg1ZYn4/MnEghhFgI
07pHgCABtpwK3RP5CDhBG/IOEsh+reztI6rd4iRcvakd4Tsaew4QWu0Rbsmo/JcI
wwMGwOE7ZtGo84Nqnk7FUA00k6jR5kSNV+cfLV00/xxunSFwZhYiY/9AQHBW9pPO
LARa/RZkm8nw7oBYYkBDOhTI/uZhApcvesX8dgNjmmdN16P40Irb/lixFu7/5g/5
YW8Elp9aqKl+KR5U1ItZf410rA/OyxzNGAn/D6PPJaiizQH42+zH/Wvks5v63hRi
J0wvdk4syhdnDxo4oKK4PU+gPduHmPwMJoSqZRQhWS5QThQM/MYvwUeOc3PKpnmh
7baFZSmK9CEIYRKrMdwzfQoZUb75FTAVWHLfFDLA0nUqiC6VKml5PlRVmrDKxb1w
37zTySz5w4Ef2PR3Nphvx5ct0SW7TW9gHQJPcRNyL9GJmvF84TkRBrwWDLj/tY34
DQeiIHJgWKnr3CSGc2/pDT4ZclCYDcy3clhMjSM/yxtWCvf7nsZisa0sVEJT70v6
tiAO126gUaffGvidl05+LCk87FELz85aqnBOW+pztOclmDIlR+AevKfVrqhS7vde

//pragma protect end_data_block
//pragma protect digest_block
2GWgggI9JtN2zqj+TElTKuljxWs=
//pragma protect end_digest_block
//pragma protect end_protected
