//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
MlpXa9nawK8v8xxKbY8Ygtuvkhm78gaGog8QRrQXJ/eT+ktjAwv35TiGZzbzO5e2
mUazlsvebCMwu8xfVbkoJAmgR1zZsMe82+opw4y7GtEZYQ5SbACkcWgPrWLL45r8
h7Q1I+AtCWzUcEUcmDPj6f6okVDzBl8hIOdIgZ5ijfk26xQ4jKi9eQ==
//pragma protect end_key_block
//pragma protect digest_block
kaKYna9xQeQ6WD3kvxh1iVsQwsc=
//pragma protect end_digest_block
//pragma protect data_block
y6TbmF8ppAl6uFrdaB84WxFkRAvQW5MWaLIkxLKULRHgxwfoPgM1RRuxYt+VU2KQ
4FBn1B2yrjMwrK6T+alGjwTaSS4GWLEK52n8E8sd+OaUsJsWZ2LexcQRF2UfGq+a
QUArLppR+U0dtb8yJt/SO2W1RQ/JsO9thldWVli0BNsOwVUXBsn4zfoMBqqb0RXe
L3lt7uicVFpuyRQUV+cR2sQuvBKF3xtx+5Px0mOTv0Y3ltG25aSSoKSlX8F5+QGF
dkTMQLik2JbNsk43KRWK602dHV+HMqRCVd8+wRx+rq/PE/le2cLbY1rUxY5nWchL
uRU0sr32R3A0t8lBMAvuuPe4FTWIfM3uTdgjGcnPCEndU0jvKeFpqjV9oaLhhEwO
u7SBg8KdeKKBV2zTiIwX+PLIptW/N+NEMoGYYwyQI65m66r61OrRx5XN0X8i6WZB
jAExDVpaWptyfOZG+JWqfk0aVxk7li8GYWiJuyq83kk1RNy1B517YAnb50VsHtu6
cmifwE3BdzYJv17z+gDAYve+XWMS5kxVNkg0qfWz+44H1p+weNrjDrn316nw20b1
0iOgXTDt8O3chFIO3IpOyJLwp7UOA0SPjdkLyqkv+gRbC1clTKqI5t14yvC6m73R
I/JpYbBwh4yiEXb/H6ViZZ0J23/KiyEh9nZfo/zEhHI08ewwB4sP/o9x7ozAl4CH
4WSyvGdtl3izyNJnzVEJb2Ez9aohm81ssrNp+gAIHU4fzhwxIGVaGJng8rvMGwzZ
yiqceYDz66bneiaPacgczqC5DQyeoZb6OWbLaMCtVvgCuglkx3KhQPhR9A0kdNeI
kqiScfamEYNS1qje5SWOjnTM0aPp6sSKMuq/7gnQ/dgIKD6o5QWETc9Kk+SWaWz4
IOC6E1BUwCbmLthUc6Ce2s++UThe4b/0xQJUBT/p+eFZ5pt0V5VRROZgDkJod1f8
rPWJ026PwJRD6YiCFhyHyxy4W9QEwOm/KwUvM4ZZ4bPQUQSSxcq/mha9AXhUwYVv
3WLnlvuSfp3SKkKvYhxs7+c41FEj6ME1x03ojclBuxXLv4W1Gh3XacQBXkpqjXxY
xtI+sHQz3jbU4RgXxzyvpQ/HgC1R9+idznwBn/xzMaUsoTbabP7zB9lML38QSUjm
EfaLCqZUdA21CzqWRRx8nCLjzYqaGSFflqJnEJknAv9gjDAA+GemrbyNZu42ezrn
udulvypDMKk9G1d14IolORxZcA/2O2RMhf9Am2hdhxFzB7uxviNJNh3JS3fMQCfS
pPL3pCo2E0Y61bPy2WHrzzT5gnOCh5wWBazuGIr0vwpfAlaXnQ46LeCZKoegarE2
h1hEObkNjICiP6UZxokT/DHCikWduku3ULXsK0hH4J7wxKLqibM2p3IidQdT/Q2R
VztT3Wj/95LqPz1DREK6mymdkgjZB7R2k3BpnSR0rGDogqIBZvax+TueT4zm/kOH
cFtvBszoN0ayuOLDiZYa16A/Q/BGj5oj9uIV1YIf3puTI9R3mCdcAIr5456IKxEX
HWV2R2uMNUTAX3B0gr2sBb13pNXLW91rMCC4RIO3BogiMqx0awILmYCeUWd1sEyN
Xyhq5ZSvZpOFhBrbClFvDL3aZZqNakW917ouPvlSI+vIx3Q/6PFlXvTJTG+n4bQK
/8zLq6U0w99b1nN7wQj3zNQ3wfzuFDKv17Ahwbb8TmTLylEGc5wbpxQrlGki96R/
cm5xCVaiWJiSfTrfXpHeUInGIkyywFE7ZSStV9H3Em9KDcTDwITknItRZ6OWEQvL
euofT6Qvw+0O/we9IiNy40mZGj0XXnSabBFRN9OSNMhTc/lkdEk43FQ2zCkZGzLV
46yqM7u2/OFzNymp8tPxWdp65Zsr9wy6o7C3rEgGDIpoFmG7gJxZm2dBS62CcTmw
+LS69uuR5pHUt+0vDsZ+lEvULpPR925ZpKJE3s+b9AMQMRXNzTvdQGwMJlymNB+5
y9N0P1O5xIZfOlp3agbNLMJrTLv4iKGQKSifmdUoiEbQqDDcdHlzNs2D/b1p2k2B
XadGD6fHQpryzUmDGYTl6hRBs8HBvmIpIVmV04jv0vx4ygzJDfggG+7z1z0ZeOii
NyQLYyGDP1MH4uc9LD77HUuMv34vX11phVipTQTDUUlIVdVhoOwq4NqZvgGRhUYq
oiduElGbOfr3ZRqSqgjp/NmXZfF9aG61/CzkP0eOtaxhayNhQN/ZjS9T3YN17A3M
TZKBuJ7tv3XFCGXCzRZOM8Tb6Y+RfZ5cuGChsS7Ph3bSAVpgheKTsvQwbntXlivN
roHkaKXk3rQ6R8OTQ9S49Z/kW76CtVfwrquZq934HG/8KmViReqZ9YzefwtVbzEc
y65DZVKPHR/SZ6fkRuAunuxGekC0W0C0d+4/qJXF5UzTT73HopIgd9mkSzkGNSd7
Mpby0t44kL+lZJoR82G6+Gd0e7OM1ggicHO65nJPuI/HkiCD6eRj/sSK05NDvGIL
UpNLB/qEcDxaO9CsAymv1Eg6unb5C9moZ0EbBjqZNfnLz00sxtH33ZPz3rrkOdSS
XNUwDcg0bRH7cVZ4VCK8lBoKSNlSfzG17HBbeUPuFXyfnlqjFjO7gGay7/9WoZQh
PbuLOcKdx9MHtDMLZumIWvJWiUMxqJrrKBerICmPO0p3cRXM/xknsdzKY/5mEs2M
gHamCJamlfAhHkDe7tkoVmwg7PFB/vG1p8mAncnA+DgJqzi2NM+zigwjg2RDJqy9
NAbkx0bNqnvKAYkGP7oechJVHcKjijhpONHfHDRptJMweBqkCsmUiuY26kLL2/U1
FMdJCDRavhsfC4/fYDvC/npuUhuALr3ZvUYUESCdZvTc7Jd07p5JjUY3htPKQaOf
NmJhZ3gLouSGXdjU3GeEcp5V4zos1v3geY3JUp3+jKtFL/XOhAZakrlefzbWM7Zb
yahRFCo54MLtjDsRPw7xDHpDlPzfvI5SLKmifoQb9OxlrFg17iRNbplwtRzjFTrL
qPlSi6w9pYWg5RRt46LL7Dp5dfDH/tXzCCugp/QMIMR7lf9a8lFnLCLv9KeR/4as
zplSC6sAQTJqt5ka/Teue6IXUlf3tPrcftuWqH7T2+OueTp+uDPk6CYJJ00Hh0sY
HOiLoUntx353TsSaGe48vetN9sNAAcXT+Rc/KXbRS0/i85AI03bXo8ei7/UURhJQ
dSsyWxj1AmLtyyAQWn346U1UvbfGsFby8tdKMxiHdc3ya7+NyqQlttBnjrfjVhTE
gzCPiOm6V1rECUAkKSak5TDqzYYfblXyr3L/HmjVy0S9VXHnbyt+OVp5LClxrgEZ
EK+HzvIk9K08/h3YZ1kL2cJdqnoe4g1vd+VZLBNHj6TRwywmSl+EVZztjnnjpx32
AJDce4qe5dFaGZVo4ov7ZVBH+kh8mItybZ0ETRjfqCa0mFfUHXXMzP74RYf21xf3
jgOWYrnmbQf/TexpthJ1z23A3IhmZra78UIGg8KQw+pVXLXv0P5Bp1j0G4hIh/ai
HTuMrGzMI5svMNjEw7fnCjsRDzmYsnN83s4HKq7k3hwQsqnoUXBAwVptbCUu2Qwz
ZkMXPvPaAbKqhZZP+Di+ClmyRxKwD7eeLnasJ2hh955zsH+8j+pi/mKL0A0jPTTo
tQHjc+TNUAbbE6Rehv/kv1/sq3ah4Fs5ql0V7OamuxTqLHgO+k51XBC+L4m5iYto
01PdEd5VmanVU8VXdeYtCT3adoIhQ6iBSUXofxhTWgbXHSaS6WwHWbsbwiAjDtTD
tkJjRa0hfgBtrWOmaHW8Zdj6boGtgCTaYG3C3HGtkimyRGES9ZgVlHgUdYDFBif3
ut7OE6c5niW3AewjNGRooSfV8al8B5Z7Py0TqmChTulQl+jJWRlfyvJ0YEzaJncS
fFoCLp45Qr3PM0wJMhIoh3xOvtbD8RpLT//PcRThi2qHd1YpUYzdybj2hXsCnGQU
6LnBP7MjD19Mw/JCoFZ2H/qZ/3S8tykg5lTkY+qnAb5uHriSUzj1uWuF3kV1RIW+
BNjzGNGfzqmHGFF0X5Nj1Te/fuGSrNUO2VkQ3/zkFri95wSLGlePoLa6oMbu7zAM
rsy0wSQzWBtoRCCoSrOHTIKHzIToVfW6+RijneSNEeCM9EfT2Z2IrQqjTgmGr+Oi
Ao9h614drG3oLqoDh5P54pYkYvJoiQL1nwbtYGoCJ0pWuHsWdJGac8+PiwKdEU6Q
wo2Twn6YHwgLn31lHQu8HrumZ/stJbP0/v/v8GtLf72AyTpMQepleRg2FdymhRXy
548339/SXKTeRSqWUKl3XFMwRYGP9byY7/l4G1T4hWn2Lgief5Vu4tIO99diGjx4
+Sv8qdObEpR0n8BgJS9b+KkUs8AbKNB5qoys8Deau5DvHpBh8TsYUBxOVIxqzZF/
LyLyBJiPrGXn/r1Ijl9EsWZCIlsMhhzKiCH30oFlp9XlQkoONBltxfAlgqRACNDH
8xN9QbA251arRw5UvnXtkbwEQzgf4SfPqLc5g3X0jOAPQ1urEqClCgD3lnkR4WgF
79vSh964uLczOuJ5n/bDwZA7EM1NOqQo6vitrJBEBcjBild6AbIqo046DasUMiB8
x+GMuYJHGB6W7mUMZcXb3s7eaXljNqdyzeMF7advALFkeyoc5LWpRcFFRo40nZMC
rC7hHYv6UvN7d4+evS5l6XSRwaJHMDKd+Fq6SK+MxX1YV4VvjeDQBmpGCMP6tAOa
GrzN0LVey2YF8YO6AYUag7oTMGTS1/ci2I5vhhDPM1soHn8TmS0KMgbh0eoJuWzs
3fQdClCfBbJ2doOFXDq3MoWbyneBRMveKmmD3hLv2P5SyPjiCgioUZ6S/vEejyzK
C+h7NEj/cF8zzllBmM6iSS0enspBzTmLwx9RxIKkJRcUMxcNUVtzFhTqSPYKDv4z
gWZWEk2NEbUnikUgFbInYGymQerauONmXl9YFibFWzY7WCHp2OBn/6Fl88DCLZPj
1dppT0UXD4ZR7+f71/MpFqCv86n8GmEZ/5LdhtjdfVZPIjHOPBqIvSRSA4zFX0xF
ryEq6ZfX7o9SdzrIpwBVijbmmHFcBUtXMLXEJy7xtizOoRwGvbIwnQqP08REzMHv
Eu0msXZ6yj739UoA4hzpFH5yfPRBqPMNAKTF7IKbD2SDFrbvxxs4yKAyRPfw5ZFs
uU3KbHs5oOmQLG2aTAdlpIMDmPuRxyc64RmGM8xNcdJqx0uyon/NLkb0/Kjx2eEM
lOpodxRDq/h440CABfesGKBBaoKCf7U/53EPCNi+qBq8oIjchVa0PaLWGjRK9CXS
ktVwgpkYaNQJDiX9dWBmGQHJ4kJDz+kY+eohYxZKa9G0KPvrMJDfiXKi7ETi7kqQ
mvLhL3aUzScyDFcVqpzlK6fBv0cDoF/R/u/JGUmHjb+H2HGvNQUefFWCdbF8S9YG
qb4PNI7l9aKfKG+5yzGF5EX3Jg0/xOb5bUiKvWV3pOnGqjpdF/a1DhO9C+pa5BqV
6/EtNo3zDU8Hx5CEWijZgkJGYvJaHYMrTNz8t4CZWSfWpa7yIrF7Y373BfPnR7k1
FiQbYAQMmtqam0DtPRL9Rj/CRgBbjyQYiwHn9Tykiwj9qaplenwpuAZ2PeWL3nIH
wlt1lEH8o5gl4LEBs1Xx7SvIenp35m2YXAj6PrCuGxTAAyTAOxTSOp7qjbhJC3n2
vbz75flHo9K4lB2f4JHdAfjoomnfimjgJHUk4njPViu3eJMH+SFydoca+ByiDAi6
gYpaJpt7Q+uprCI+6GyNoEurjx5kdOZx0gSb3JryloEMhyRw63FAaPkMMbLg0SzJ
GOiAyh0lj1qidrQPCo6c4/sA7IwbcmGLMPvRsCv2ogNGV8BjOv28c6Pb7MW7IEHo
+S5zIDMrBt95NJCXtHUyStGbFJZ3xPYndsfg80NG7fut3SlV8Cdww8k+JYXv39Ef
cI7h1k6PMn7RtPGRCR45A272GCvknU+2ZBXQ+zR6/tAQQrHbLHlFhkoXSrSzK53y
NtflyFNI9Jv06XIgKYNMbUhcraQTPVbGA5OkcMlUDrksgZnsj2l6wmIxwGzbl1Vd
a2qbO+qbS3TPqs28gQ/P341lOr1WvO/W107dnAtz+ul3D9K8av96x9fXvjkG7lEp
AC5QWlzgGohPULl77/s+E5/2ghCWJdVuKMyWEMbfd23xe1+XvCPBN1GwjQ+QyWii
c9LSX+XWyGJZOjsAOjfivNyJTpM2gnlKfUVViNsKI4DspiSlzkTRq+IoOhqEemz0
LRQiEOa5OTh5Gh/hHiJtsTS4vzv0wK0mFy41hag/ML6lAS5t6L3UxZTZzjPx+fwf
aYAnxhf1+dTbm1vl6P48uSCbWf1PmkPcqwngUN53DxF8jX4Ah7D/dMkWnQ381bUl
9aka3FIaOL6XVn5MHv7bd19r3kZQiSytdzJNgj1YuSpq7NarRAB6utc+ScO2oT5n
7tRBKCJ2GzZGb+yMoa/pO1e6VhEUoUNiuom+ZEzuhuw4XZXjaSwv/TmOnWnNBFdC
3l96R3uhzS/Z6vaMegJOYgNdj9xYbUfe5EON2FTCdgGKWj1sK2fPI+iG98hCP8rJ
giV46q+yMxBwuBcmnZNGKka0e6awWDjEmdjrW4Ni2/17rXXd0BxTK5McqkGA+nfU
r1sQXYtvCKK9lPkXpDF9oqe7UXrp3OqMEBmdEdTkBY8GJ/+1Id803TCIf2YlQpXf
RAVlxJ9vGOfNwdhcsnc+a7FPQTdffLRoQaB5f0fvQxmCuCTdG/NHnxzbkEszP8Jd
TFpRUdV2LBMQH/uupz7R1f/67DW64Or0SwtU/PDDiu2k15EBzL5uXrbtiXFfof0k
RWIKnVNr0Rq6WKXne4mfcG0xw7p2eklFmzyLuFyTU/ieEmqBhOkGI5Lk+sz9wKDE
BkRkvOXqtMJeVS/Gg7jy9f4UmMWGTRdGYgB90SKCk9ZbIMkfCs2r5BnzS3mJNVI3
36Z5JDW6udqaZKESr4R2eIRsXMg1p/39xnovCqmz36LTSOGOE0Ha+KiSU9Fb0eKW
FPlW0OYMio3blBsxOiBBxm2LtB5GYmwIohvERAl2vgdZSkjsMr+831jYAWGLQT4b
Bf056S8iRivyXi5AYEJKDKNUZlRikhI/T+oZjL3gTfCxx8caZywIdPoMa7ppP//z
iJtbwhLDA88J7Xpi23YWGkH7d2T7E7pIlctUiJbiJxiozgyenbakGbzFnLQRACyr
KocOzBHJmCfzftORd0GhRvQyjze7T1yJq7UzjVKZd14xUlhJ2e5IFXfPGMjI1gaj
kQ+1eq9AG3URscHwFfQNh4YR6ivYyhddk+i+eGjNyw8DPjqqkHkKI/K8JN3IaAYa
0JK3GO1lcSPdrdLCMAC5oIUMWf0EpTEuBlKY9xqH2HN1zG6JPtlXmcjSGUdTFK41
wWe5ZnVk+XZYUgqKu7WMIqTdKLXNO3q6hN2Wlue8M7LyjuBIaOPi/TbWE3v6NBOD
o0UEsUWu31ykyDw7s25IMXOblHckcH/xAXITpr7FWyS6FDdKo/s1ClxCeh1DpzuE
Bosamfj51kLlED3HC3QpdkE7snCdMwGhQGpqx879ZBuQBnRnzFtNPQnD2oinrn6Y
F5uuKTsSui4NFHTiDiuOaLcctSp3xU9Wk2wcDx6w7rO2FQutHRrep4VTSKmNT+np
1Gqqp7Hf1DCcCgvOd42gjEJ2OvSxnvliJjs5dKhvE9SHpFtrONVn8ySYs302bHnF
i89/24W7jzaga7k2kh+aPVBYyUR9uMfN3X9apQ+Lc9SK1uoHFMgK6BoAEkN3i3sF
dXd1h8fCBaQ9jPLq3tOmHulLxIgxpK8oe+WurlB17d7vJohPQW6J0PoFrq0Vrd22
eRAtgAOjyK/nk9fIknC34REUNPvmlB8wrPtELkCSVivCLDN1iTR7OJmEoq6JQHfk
2WIRiJwlcqoMeanXw8MfNNn20IXXc2JkTiwHsQNi3RKfX/1tqlgeeTi7Mvzt7Y7T
kOh9Z9CI58ePAwMEt2R2M1VmRwIKj2k33u6jywAKvAJWtDJo3IbPpaVzowr09Ch/
dk43+dAXcMANhRCSy5vHIc00czL6/MTTcaeunCyttAg29ZC8X6090kw0kFxCFoWH
0lnhumoNrFcrKDxEbabFpiCzeYVwvAqajnnGufVaZk3AZoWcLY+faWKjmXlZ3haj
5AjADPog17iJbZdaPNPRn3b+eWjz9jSGTEzhll6MHJw5YyTNkB4ekWwQ+pdC68K/
2MTLhlhAuwKTuJjmXeb2opBabP5agpby0mTfzuPhkaPc2J1Dj0vQ8czk3MOSIo3X
UifEpDzwR9atAuJ1LaA8MQNo6Qz8MI5C28uKH3p+VI331648FjN8I9FZrSQ8IEpM
EZQcBulYY5dXZKt9qLP+10QDf0tPptUFwod6wY5qegCSPTAM0sgyJM/PRI70a7Lr
Jr3PGzR3K9En/61nOnrvd0g0ke+PZAlczB37GAmtSjHw/LbZ5elBzF4uSf537Cpe
fJptji9zRkLKQI99oVw8gjyJim8zT8dPHbQajedTcnxBX9/vcHGYXjXIG4vaCKD7
5pbnrBxmeNoxmTwLrIEe7LQx0hVzvVJcSce+znlavU3XR4WHxqq0QAoOcUA2Bqiq
+hexAd5EUpsFjwSPGV4YHn5O2EiaCV5xVn7a1pO8T++kZ6o6a7X4ihTgK4IVIxk8
+KISX4GEX42EV/Hj+b9DYVTPovzcpRhQQee8Ih3rVoXvyPJ1NcbE7l/q7YxwEGmT
S/YqVOwez95Jys8HUz88MF1YKEgrZzKbXrE20UiibBdqAaQZRuT6HqWcMA/O4Ixx
6a7e2i+tn5e03qldFUMBZK3FDjTIU7BCkDnbynVPXDxhY33hL1Y67LHTF0vDGyrA
EewHZlh55wFNKzmvee6nKN6Kw6IFNKQsvBQw8XGwwp/0zyDw5j8oPazcaM7z1LdW
9/e9S+5eWrJHOLhWF30GEOnWAGUTAuVEmf2JoVsBZiKB2HwGwUVAwNkBEfgYoMlP
1kuMt2OeC9A6UjrcV/Gap0reb1rbAGbx41H/vfBBttQsJ7rlMKjYVFF8fgM+/254
37SxgYxbgC9syvosOaJ1efgtzweQ/+QskiWprTQaCXfbdUqAoXsTK65RfHKY5ZMT
TY1R4RR1BbtWTENikPviMT8kXinp7+O3FqoeOPhumgamW55EsXnntFdMQkQs8RQK
FsQsseOhRn948Xv6cE4Gsyjoe2lc6E2CqIpwy2oOVc7vbyMw2mETG3oo7b39Gegj
3Y/NLNtsWGjpnhg6IljhFvMe97sj5FpHnOhvy5uNoUurhxfZ+Lz23/j1BH7xAYHZ
UckNTewdQm61P6S/SMn78s96tkTdJqFq698vSwfOteFvVlcfoJh1nTJT5qab0Lo0
pUztY6wkbhExj5PaZetTER1FuuuAC/tF4KN63uS51J43L3vAOmhBjmxi+sPiCzs1
4mcjR66F6/Cq+fBMAXB9k/pJkHwmnk47q6alVBzVmgBMuBsmC6HGwpkaqa1sfr9V
+wk1XP+4oh9s6ZYmpXrc89CoH27fhCailhk1JMqqgDdeRcxotgHNn/KAYnGyg8TR
rbo5bsjD3zD30HXjjkzAihmci5yUiCKe1zeJLXprCag/ddAhqfAfYQ93qlS3xG0/
McG7s+14bD1MUbWKJVQS9RqrU80AdTzLJe8SwDkXfWi5RNcL9P6kwXoBo+nA+BAP
naEQuxzQP5Z/OZKKIUMxbR5yzloH+q+ivcjhVvSV1QVgNp9eev9bsCRnn7/+r+3P
KnFv7NMEKgFXoN+5hXFkYBQ0exVVZCMe5MQ/+xSAXlA2WX2fADroBOtOjCGCzyK2
tKfYKj6gUFr148zhifx6stiul44ivBNa/ixTFqQy4q4BidAP+CWD9q8GqAmq4ivX
vP8o8Z0HJGCyiZf/LFifit+ndOGR0XtnjE86wUruY5UzeBxls85thUbLqpRS+TqA
j6OSn+VLtf0QMVcFgVX9kdWWwJf5+OYzI7miWjjbyde8wXlYB3wCdHce2mpVP8D2
oTr6PSGEqOS+YZmEqG2XevZEUyvm0YrqZJiJrzeEC8so2ughgPepQHAAUguKsOgM
hLb3ctK83xqhBqIxHFenDTjQKO5uPTAHhxPhqiorRYgSOWgSKHxq1O1vm6PPQA7H
YmaLO663oqM9UelquuMhRc9p67ToX1jX7qV5enA7Jm7eKpVA4aOg2My/bV/VsOQr
5uCeVAXxD0Y8QtjYLy9IwlJisisQhaBDpqamf1H5knj5CeplLoA6djtAb1LXsCb+
Tnq/exzj8XgTLwACH3O7vo5JWkhFj38fLjnruiwAuewGzHNS+HcnuP+7kByyqlvD
JTXWEeSJ3Jxp4QfGyFWD1fNm09SqRlKcrws0l0X+0pUETabes3H3nJliV0vU2hmF
lDJe/Q+bZFG9UkD3TUlQUaiwTyWABa0DUBeTb0ClGniiKQrj7bZ5qfrGq2Xwioj7
Lh8aHo/PWGwBiLwxWdYwJy5skpV5ii7/IsGUsOO98DT7eAAmXuZvlsAcW69Fe6NE
fPBeGRlPiEgJuxcX7yLrbK0Cq7/74A9oP2gaKXIlVZVRVgQYmdNCA1k3jI2UZjZk
sydZcsPxDuXlLXCMRlVrSLbjSBr2LAK1jzqQxKzV8rEToyQ3s+p4xx3tTqOHbvD4
kzdre2axS9Il6gmIU/vlD+hY6POoD1icMHYJCEsS9G99tkBWITv10k8RQNYdm3pe
xZ6D1HeBB3rGdknIuU6J9L78R8IhNC+ND3wwLltGfCRqfRd6TFqNGpxBXsA5GVSd
JKicBmEF4J6+Kj+pBAa27pGbQDmIJQ9MIuE0+ez7yF6zujEke1GsldqxvS2Suvbw
GYgtsHKgHBKI+zIPLQBG7Kma7tZvI7V/5wLrxcIeXecmQb4qJkJtzAEoRLPbsRgU
YoeGPIbVukdeV54w3dL5B0P/eS0sbMiuEN8dnyADHB43pSzRavg0Y/rlWL7ip3fX
GMQiQPyoKfjOZz1eAQ+oTZgJTIZojYKMNw/kQRFq1lOLXOmw9SaX63eg5IdIZK6f
siY/hdY4OB3wnlmRUsTughYz27nWMJ0t3+sJmclCeQvmdhWbPTYUrutkh7Lmp1tz
tzUHAUjEjrfIK3ReQJ7Jl3Vvk+K+x3qfh1xiGhHtNFGeWIa5Q07hpO83h7Z6DTKc
l2StkUvjVrCw0ftv9h1IOXAlbZSyI5u2zs0d8u6LSDtjXDKF/fNNsejCM/sRvw2j
kKyEJ2DSFG/Pg5Vs0K4gDj8wrsZrf9cWNT/XEBUzsQHR7OFK+sVLp2tk4+YMkx3+
bfRToJjKRazSUkj1pFOowbIfAgi7JYDCGspbejkN/YmU7CDyv/2O1jMliQbsC2R9
DyUYXT/5H0nOGI/X88skjDOennooAnG7SbssilO7pYs+Nvl/Of9rY1zAtGOONyTS
p9oI8ZmyAH9hrlAD0tRyVCE63Z/WSXOiJonfCIqLYlgpICuli4gPa4kTlLQ2vvy1
PXT3AqpXHC/9smwzMZjkt/WQxISX4YXIuwSKESe9tHeNv02pnwvFWpg0sfKJwz7Z
Y2fhqIwEYEv3Fl27oljomOoLwGaZlDM0Ui+eASN2UjaQf4nUKMM66plND9p8a4CD
91tHj2+UMt1hWpMCU2KUwYeECNMUL2NDKFtazT7EMH4wLKGv/W2XpFMcCxSdm8Hz
5gWmsIJOVg2m8zDAlTrfs4vvjk+nCwGGqOkeuXZA8Me/jJyTPuLCAczpstdF+Ugy
7I6yeh95j+VQG0CI0tzIdb6E9nKoVndWFHbpc9RSm+kgHYMdXTjN2z0d9/NWnx+A
DzxsFBfNBvZD8R9Y6ZI34S6Utk3iLR9sXH9WL3y+BPRso1lNwr+nIc5PX0/0KJT/
QauXqN3An3XNlzlGS1YcsQlouQ8HYjEoCudD88CxnhKPLkFx/8lw9zsyK0cTS+Wh
wGYXnzxqNXIG5stcEIv+nDiEnWSwumaT2h/DwZeGHJtajwOcwprLOf2xP06SES3h
/z7a7+8cuOnEA7p4iNuk7jUDAiqX/2oDxmJMVCCLG4rDupvseGF3rZVXSwkP22Lr
DH8+3BoWwg7nGieMC1W67hH+Hg6cWCQv2ISXbSL78VKiQYejmOQVwXWf6e5Pg5eH
N0d2wrI7/NlMiOberZGc4Po/uyTi6jjkBmlSfY5QxuBSyTu9boBWLPnZFmFEFjUX
z/zswBbNutuXz024DTzj+EeBliMgVICZRoPT5tKhXwXnHUsIsgcEjNF1/3GuzlO1
m2bOyMJkoI1O2PaA6cxvZHEdz49xYFcemKsR3gBLtkMqaxBQBTYnbHA2O5N2yjJb
/tMQsmEK9lD+91ZK45pSp8jodUP9YCT6vfS83kJgss7FvlQzTV5EncN5Jb51iJcO
xIfynYrH4Wlw9FUcvfwWsEYlE7RxLRgxFAImdDmVrI5W9cgncHpnsSvPSru6RppN
C/vFFxqAAtXJbueIehWTcpewOjvPncBaCBfBsKMvskwSz/oGTehYNVy34VEavTLG
UyOobA/658YG/Oa+ZgplGgquFgBnuJFzxjnnsqzzrWMKm2TYIlmAVvFnIL/gcXpo
BwQYrnhjOcBK7jirWEiyL8lUQ1YrRZaKwkgb8jge76V8cAtcesqm5jeKBZrpVCjt
st+j+UMGqbXsrcstzQEBXJjQt+TpwaSItp+IHworPiSz91FbHu++MT6TyQhg3Sf8
wO8xyMmUo5nH4q6JMYFMxpTsA9tkckVrhVKl94Q+er3kfMB+ShmwwCNJ5ULRUJNa
NB7MUFD+jLT8N4I+nyk8qOtxArn+hPCkSmJ9E1D9NJZYr69leCIqoZ7AfNx+Xj9i
J49TrtTe6K6iqK9ksYZR9ttHRZH2YArsB+MP6TpNUHpM7QU/Zxi4yFqzAWCjb+2D
XjD4rsBzYpeVdx0fnFomDA6uquweK7/VDWRTUzymmOt0TFq+ujOol3/EGPNR6Khi
NT8z31HE9S88WAInshiDdUDYjtXIDusVKEyHQrUS48xMPcLw+M8WQEFp3/eldcdk
dFXAo+BkZJ/rWYCAhXlRaY/f7TD0Om84ekCGmgC5btsjlN2iHZMC29OEk3xyV/8d
2YeHrmW20zSd6+5ztEFQSGErUbbGlksAewHvJQWUrqSiMFI/CmdnZli6APHUGhdh
Fpk4MZt0EyH5zVRDVJun8ruMEUlR12n+rDmYO1NO1emGlnGrXI5/Vylops0chzuP
RVz6QsUkwzdYFlJ0ZbO8I4VcTqX2AxcsXCaJZQY9jmWcCA+q+/TeHkR/Vrh3FJ/Q
P0Zc1HnW7sj9qWeH87X26rVjDz45c1CiWslk+LdscEbL0hmOUgd6Si1uK5AeyeaA
hAsgeTn62sIFCqV8nVUQCNvWtIJAz4qBk28xGMQoloyLiEFWp/D/7k65LkKEIqpi
8PMiyJF/fOxDat7KVHhbIMIt3BGrTWJYhxNInIqOST6pOw+HMjhb9qNO0vnGlSAD
eAjtBeA8SSV4G9QdoOpOGH39I5w65pjBSkY/ojGkv84czhzexrGR52UNdA/ZOAt9
Ede4GKyjbNbLojY2eyM/RkbfjNyaXl57IHNqOjmtvkKC35f9qLiOz6ZsEUre7NpN
kQZlKvZfIwa2/vzsXpAz1aB+wJXitzNcA3RURWcmXarsY30ODbFMKlyaCj1wBCdL
Ej158O0v0V2HfGICiVb5nn56fhjF8Eh07LP0XQsGBeXyYv7QXNjRI8cuS7dL4NOU
jJk6itLDZ0t5+E+BsN3uTbOpUddPtkl4VhozWy8dfONvNQsqmVXGjW9qGE7Geeec
CI/B9FqBQKiiU/SahrqwGM5OWMdOB0g7F9M/P5eq1i0RcnLvMafMH5+UwUW+o6E7
9R+/A9ALvHO0nNCmGgp8yzNT+GbQ3V9/eVEMe9I/X3NOmIPs91O4YWf79EExi4ks
Rl9mZMotKOW0e7xLrxZ9vnedg/lo0s1zOex4kIfHXuGWOeC/xpZnr7RHXRsej0Vg
UpXeOjroLL1aeFFEyJ4XhMb0usecNo4jcMCtDpPMlxv9/buO3lLNlWtPJgtOofno
bk5TLUSUSKZ5m/JC4TBJeMC3Wc8ysfYh8t5oVb3up50L2yZ6egdwuFW9JEwwBr1+
eRpDgeQOvFhTEmzUQZnGuhu7+sjgVSil+ZKQz2DxNoqAKK8E+NbfSh0zrwAaeOAE
bXZQ7EKDhFnHJDuCDvoEe8dpMQNn6Vym/2MJ/YptK0zdsrqgpaWpGc0Tpo8Vebqy
Uqm0oaLXlc4/1jrAteatqNhQJ4y5Bl1P+oTYES6l5dtIn4nnTUmUNnHtm2LejwbC
jxW1c51wXzaY0KZ3Q3JugicUWUwMuFayUQnuWaR8LSSjJtBB70JtiEKudt53r34D
aoXE+yvQazd9yCG+jfQ/R+hLevMkW+nf9OIbcDl/sMB5CCBBz9/kkUV7IxqTgBL0
D4hXe1IrKaYxGegqjhCkMuG21xJEQV8wKWWEQfuYaZtxFfvtlEu+mt422yxvCc+O
grjoUJYvL53Wmn4gO8guC7ogcaeIopH8pEHHq8ZYQPYd/cpjZFEvBocmfHRoEp0U
QvTDBmmF1ZZUtNAJ8WnD78ayf0Sl4SDAohnL7rWuqlTYNWQVzLJf3UDzyBs2M82K
BGfimmusdkmUuNMUt2pbzupas1l7emS15trZEZuCiJelAnacRBscs/324KquSI8K
uVQDecqcPIcX5do8Rxv54Q6EEBI8vk/fYazokdFa3m7oEVNS4Ez2LUlG4JMI/esC
GcTRVro6nLT7Po3yNweBb+AiD8NrfFpqiB/UKlp6ZjMv0gw3NLbWFnktqJV+BZNc
rakR3FT/hTf7bmqIpIr7n8GiHMd82OYlvPQhbEh3wRjbvDX1Da1YE94hrYOXKyTi
MOf68xfqb4wMN7qjssgYwMT5DSnFm320yG2dWAFnpnCmgXRnh61VN3pu7cC5zPHy
Rj37+x6CI/+RpnDq5a4vzkc2qs/f0STfXKEaWKZGiJn9wBPgPhoEQIr/UQCMsN8g
GE7LFk66MG+DUIHDKYd00DhWn1LVoJKUE29EFGvuBz+zCBWmZtrUwKM1bhZ+NRHM
+GLn6J9Ta/sSJOaAnc0z8EsXOC3cUww7Us5fpG9bJBSIDjSmPfXYKPOHdZJ+2EgQ
aZKKsQN6JLbTUQ3xPsiQ0u4wi1W4xCLHgvipzGALQvjBCHcTy190SydfOK+z0g3/
895T/Zvhh66zGzysyjaFhR6zhOPL1BTTBQ/JHlJAajF8Ug+Vf4MDrsF+g3r26FEC
BtiPvxeWCLlEawWlCPmUjVYwpPtkDE3uH6ogZ4ziR4dCEk0N8zwIjDHJ/CPO4V4j
ElrMNRx92MTNUgqeMp+2WjR+T3tdUnLErElbW/fvSJR083nQAH7nJr8fT7tOVYNy
ZjN4BuBxprHFrBFRKdkJuXpBrM1dtQAIPpoP3QwrXInqJwdcm2TjvwRnqxPG3dDp
9jFwf9floJtD6MYSJusaGGj+S+0KsCOSInKF0xeZY+ZowdKYmvbXi5dBid8Fzhdb
Sw/sHfFegOlGhaGKy5NScKf9HcfvFOklZD+Ht7+1r5T5RY8/ovyWOAIbL4BgDsAC
aK5c1/vd5qBgvye9LGuxj/BYvoEvmbftaAKzdTlpZsCA7CcJvahYdLoEA+37o+2W
EqiWmQGfGusr5yLBAL4YH1yPpDLRC2P+WH26xKqprRQn54gi1JkEKfxT/N6X5HXd
+lWKnlEq52iqQaWYyBkmgzbckQuz4JmN2re81pgBcMM/s6V35GvwjWb2fSmRJwN9
DyxbYXC4P84j61pgszDfUEg/tcnQXktCUAI8TjryTfZp1xP2OabmIuXActTg+lZy
f0gWPDWDX8Jdbf3TvN94rGxWXs6LwpLyi3pKgZFSSiNXz+f4xeAaqHqUlUEEji6i
NDisjdH/c1pSnhstrWmGj3EIK/67nqIk3Id0FiG1IprFcJhu1l8iQcL7XjU/96U6
MveV2vGEgONxr3n3vRQ55w9AD8g/mp5u6iOv0/Z3Q1GawuT8ltOf4jSn8R18zifI
7Aq+c2HgSd5jwS/r7BzQLMIhSmyoRryJgx73Ntcd//QmDdFoHTwhQCghOye5xCGH
Yum81zZnraUYf/nR+/xNP9pEqpVM401XAn+4t96PA4ud7xKH5Hv7mrmlx6Y4ArRD
ocDj5IzTOekc11Pa+6Q4vwUNXF3QH3KwAZBOexwlP/ZVZP+j1tgZZgu9HdQpBMmS
H9WtEmXr1mivxDVyUscgYwu3ngzUQB+TDZ4UJQEBPJrjQpp2r9lvswIDIrnm6qQS
1EMzGhbJ5j0HXagzVi1RF3+fsOM59gMUGoG5SAyoZRMySbCVSE2hZY9HfQi/13fD
+Y5KiOXbP1EXNwVk2vBXVUwFqOGzWk/B6HCLMuD7gNmi2Dx/bFI8j4/h1q+P84jS
vKkhbyV9mkPT5oOTWe6qvQA6D6nO6MD+cqKHtDHYPVazzY7Iw9HNBFhENjv49UGv
gQhOmmIkc9PUOsmGj78k9CgXPzTdLGyxOz72thvuQ5f3QzepbdVzjfWiteEshsNa
8PVHCxmAj/dTQa35SWoftfpjV36FU36Fyf0joZqJWvKO1WSwM68w+9GEJs+z6OKh
C28llgzCvmGnHbAJsVu4E5frSuO/DKU1F1T3oSASMqiR7r5EYuLSURA/botQ/MUN
l54kmgpwO8WolqLW6twkKiQu8ffjYAMj7ZK3adqtSvHUzSCYDJZGwq+2Uyq8g7iH
/DoGGmnXR+RdDIauaoLMXveYE8dSd6O0Uyd22URszHTNN4gjzrPXr1b75K2rGAPx
Ii0+QUoH3oW4upwLCyOx3ogxR7PI0iJyii0YyUsTUxSqLFtPVoLhxWtbLy/x3QSv
1saN4aY+1OHGq/2kac4hEgopKukByGJ5XFkl/qy/1EfFG2OD55ybu74K4tQBO/te
/9reNjulBbh3lUeZf4rKvtfS4B+HpcWPDy+xy8Tl4WaVMPTz8W9GN0t+Gdyezvbe
JMhFcCA7AxM4KmDoP/t7ujJzQlLiUpLIy1kSJESfgijzPPlIejy0lPesTbnpgoRz
DdteEvvvf3XRUeTUSw/vG2zTOskUV2eDFk+c8hmEoIsCVJ4uB0OKcwTpHEzcKQvD
pP/LacIrTCA8lBwX4/k1osbkh8quHq/XQubnQR1VgzwPGjD80AbNIy9JCZpJ1j58
R/6dfxirHffQ6ENLA5skF4rGLOU2+Oeo7cqDtBZaS0XscsitZsvszVWJWTxy5FY1
BJJlbunugFAiyY5k7CT7Gr4bXdhCG/kl+fRZk9cH4wvVkOdU8mxVW7s3wEBDcHFZ
yZH1YX26SY5C4y7NmCX2T/7n+bkD9OwwQFt0vf8HfmNSdKRbaA6kr0q0CzLE8gk+
r1Hdjgo6Xs07WrEUbk7xcc+OEfTsr7Yn6pS4OomQ3uBPP9KTJn5PF93IcxW0mdey
0/FCcpNxgCwOpFQ6s07DKsWrx5xn1qv+4I0LQRpbwc9kNCym+tWVXacJkO19BF6c
cux/FN/cgNX4e2O/qFTn5qzPBi9155AUTR2bfYlpRGcMu/CuZgCxG636lw9eZuOi
IbTp4MDwbRnbNuchJkWAEu2fqK3AkEmU5NZ+e3hMd7AMvRMgCDylyjDZqWBu0v/V
e9izappnZZZjADmgfLz9ZE9jc9OGGsAHayR2vrU5gkhxRMd8AxmCiiK9CFSvXOqN
Zbo+ojiGLaDr7gB/yrTDeZKeYsIivWYhNcUQG5M54F62Ksk6o+dCvVUJEDylTatQ
snRswHNysGS7BnVaUMljkRVMdrnrXkNjK4SEzI1FQH8h3wagNCuAwELyT6irDDQp
98dZRSO4SLRfet+UFVJe0QbgMUUafYUa+UpYV4auxG7aIXKROpdJ8C/I+gfp+HLx
HcUGde3/pngoZ5aNJxbILsxCpVSX6Z0fakSVB5NgWOjM5D65XfTECMHac8xvBMVk
B+NWyo8m/Xwouu+1b0Ki7JI9hU5DHk0xc35X9Bf9moUFF18FW5eQYLDc2oBc3/cR
LYiwvrL9Ny58xwemZqoXpTkInI2gUDcmCtRQxVOuDnQ6CMHCFpH3ldeHOpCxkAER
A5Nc6pO03XURMNig+km90AuiH2soxu/lKrLLIY4geQ5iX5Y/uwIQOnP27k+uZbva
APyhP8gSd7mFNa3QEwZcU2H8jjrwLZ1Yf95ETDO0Gv/Cw1eZGvIpsu4un5u3wF1f
W0lZvst2PyNHUdnljp2EL8uP+IV9UFISGnSxvL7sqzHuBEFxIPHaQ7PgkiEyYP2C
7coDAJmJUQBpKNoeMcXaxix08o0r68/xYfbDq4lYz+VSMIERV04gv1yJnlR6DdhG
KRKxJK3lxJDHLbziSr6ePOHyGAcOm+BuhVqzDrvtdAX3VslEqrq2clqJnJ3aIrSO
tbNnYtdBRZnVDx1dNLw3Gld+jaEUss/cFiI1MawROTEtEECL5YGCqRdopdXYTMfC
Bv5vIuIaykhfJa2/2gm0DC25rjhM4/ZCU5ah3TRs/cX9gVSE9XmFMjX/knI4YfYl
YBYcgUCA6j6RWWogN5jFV4MwX1zMa7jGao8SEBlswsBj8I4AP7AdiN2jdh8zAXNr
WrplGRHbWWne1cKpiljDnFSq40Rn6g76OZ/HttUOfedKB4dng0DC5oNPyQK5XJLc
DzYDWhGzDBMPYY2ofoGTcm2eJXEHK8CtApW/fF/Lfd5Hf4x/u6TC8f2GYTJe+hX2
Wcm91RDooWuwI5W77NAFaDXdGr51STuoak4NlHlkRT4gSv/NZuReD/x9a4yGuajc
enc5nH6g3wdIJPytw0hmszI+YOfkNhoneDZKc+woM4lg0b9BfISdPhdKnLD9kJwv
BrrXSr2dIjDltYEG4AV2ibjdK6Li3uLZR5hnTS2df+DRn5i5t8Im3Srm8r1F52DO
YG7mSHkGCf8RFjuc1I4syCpL0UsEmbQkslpm4eQxs4c2iEzas/uE1btHE6INvC6e
YbknHkqU3LHT7kVAeHPVnDpA/x6m5C6TMaXE1bSn3XP9sPYyqIwQSav0edQ6YGkr
B2+mVmw183JrGkG1FY8hbYKwUNUnhQvtd3nuUJjdLOXX+jAZiPQowbhqlQcWwqj4
yYWZL1MsFxswiNxU+r5J1y9epL1+ijBNA7OjsZ+o1Bs7Ij1UpOSKr5prXXj2ed9n
3VE7pH1k+DdDQRvDT2dO5KyuNCbmGB/892Y8Tf5Ira028+aITInQEx4JGJF03/NU
dn4rlRC1AQgqL1HVNe3n9MzHFsQEaFkgdIXXe3XLXqMmqsu7y1cY5rXZCXA1cIHu
oLWO1VeFGznd3gSjMYdoYeBxzQbNhzQJqWjhs73+O9qp61LK/OvumoPSpugeEJvk
QyYlc8Zt3f9si/WNVunsNQwUttOqxtY3qhki14O0Nda6C8kGPmz8QpAXQ66wpL/k
rTqYS9TrrWiUc+7cdlsCyDV03P71oxyKnUqzvewum3khicAnBQP+NTZf9MN7GoUL
tukTXdDxrJivP0e+as21t2mHZKb73HkHiGp+kaAfDIzlZB4pq8OFBlLRlt7cDqFL
qmouPJBZ3hUebXlotpMj84UtaRqG+eM0xi+in34jf2o9MVoKebvtJ0/f76jqqrfi
T/HUwvA3Ug3SJPsox5+Nq5XSpuK1ExRT56fN39xke8xTjY5Gmb2f2RqghihSv261
h+gDu4/jqk1bUomHBVVqQV1PLfIUvJ5al0Gg8O8RkKEU3B5kccndYDLq1XCnk7+B
0Pa2eG3peNVZjTwAGmT/H6TasyQyLsTKJaNe0tWCD7HgaqSK70l9LVU7oN1cge7z
OFZM80EDoRx5ThdUcTtGKs+Wjz+DKALLnmqJbCQQ+ofQw5apL9qh9pBukXvnzpeh
FLCNjrDXQki9/CdIERZAaR8UXUpV4ezQBsAPi0pSWbBb6Xgnp8Ye8Hse484Q+Hsx
qEVEvsCKeN0s/+9svbAEfUAT2FHs0LauuPtLAOp37Tg6TosQxop2DrL5mbJzNx0i
HJc1WXuA7nHcnpcO/49P9WExt9Oe6aehPL75JeNcG/aaA9Vb3GphrDl0rJUDgKQZ
An5AjJn3H14wz9SRvrqdW1fKsQOK6U1XYjQoGoIYyO67Nz/X5eqq085/pQzmkdpT
N3rJVHr5ounHzqz7+FQM5D8vUlebYOCayXKGaw6wjl2a+0zfxg35AjfpGPNlBbjJ
9etj7BnpkMd7ci4y4j16L9TNWRntDdTDLdTPMdre1NCsF0nwkZ8Hqr2QGu0ue1n/
Yhk/+TIvOXW9fqAQbnRU3WUVGJS2eECSmNOUIVLx+7heddv2x4XUi/C9FrRmUTUe
a2fKMz3x1TmfliPLBlPQjHyoolzv+Rj4jzbFfycr3RuAVfQBfLuPdet/G2jFq4yz
qP+N7Q+2iEn6uSxdzk/gDHMwYoT0UvcIxlvvRGgSwwEatKoSG9AUwa27j+dv/2TE
LBeFm55bpQhpoFKZpE0SpaEwJwAOuwvL1+9gAvx9Uw4lZQPNW0GfB0FOiJWr+wNX
A1j7OjJ9UV0AMIqqNqH6+GDOGXCDZvqLKuZ1/qLowzDDNhyX/d8ZrNizScBc+PVI
Xp+WbcYeNzOQZzA4NbA0dBpObHoWtjx+GBcE6KR8KewdUxmvBkaAktfK9LfwNc4x
JLJMPWSVChLEZYSInnVVeQHdy1ueQ4sk5TK46UpQqkmWnhScFn1Y3f8YgnBuLaIK
Q3Xngqf9ITeQBb3aaemzA+FjMxkJuWUBSb+IVtH9gkJGs+rqymD35AjZqIs0j6yM
c7RJxsV/MlfcF79xpuHWkrmTJxhlPG+sni0HAS1m2MIV78KVCOjYZe6ZrOqRwkdf
6bu/9IBAJPMf+TMfR7zA9i/nQALaMcWrGLHRuCoaLHGYDgQ7jzDiqnZf+O3jLxdF
ZfWZ6/AlhInKxc/+RGW6sR7n9NY27vKSqMdxX3bt7/uGbTqF4/Popt+3m05ymME3
QOkEJNhBMuvbeOryY2ojJIXU5FxYK4jeRLUg/3AKdi3pXWIf5YLAAD+M1eYAvr+W
nF+wKy5rcK0tZUaGOlRUbbN2ZOtzNGfYS7j76eZq1Y35MEV8hJdSxLW24dCtFZhO
Jp8IoIYP0l0O9mCWCpz5tS5z4dOI77MwHf5ANjCu2BHrCCWE/phM4svEXefQ2aKL
Whu2pTXFyQzawvFyG++bj39KvggAayIMMUrW6UC+zh9I9QIp+yEOWis8rznSJnGZ
yZ4sECX/t7fBH3dvqH7xPuuHrLLCyQtZjM7EKaCXH2q6kkHs7xx9w3ZzFxn+z6qt
+zUFr4kyDJTzOIxlgpnsQ6kkS02/mylQL82RXdZvECX6AXWkc+VYk+D/YAIIUHQK
bqEsOIcl8UaRkF/GCiZJ1uMVBh1Vc1SE7Lr7pfq5phrRYn6kuevacWwXLkuk2PvT
M/k82KOJ7KR4nrUnhuTnzm+iSiI6l5+UjFzOnBQWWh98gJvKgya+q8sATxiMUj18
sZCmChoi1zpk0SUXJYqLaxIO5aG/5fusQ/xEUcBagyt6f2OMNJ2maVeqlACzC86M
TjEv98foInxSWozXBte2YILN2BHHaf9dvR0OmNklK+gXifFNGT0/y+T2gv303QHY
KsyvdpL/T+Lq97oDI/VmdDzWW3HrAimLaSY/lV9j7FhUK+iEuQPJDvkmfl18CWCX
DbfnyaNCIwJGeUALv9H0E2p2bHSgoMHrFB4JM4woqyNaIA36ilVA6TYcj3Ck0Yr8
rtXiCLqPEvvHqR2jwr2IDM71Ie0WJcoxASveA7GmbcUCreQ/j+z9iEhlv5FDpa1T
Y2j5ULvg5v2FmdkdXSvL8FsmMW51XguciX2CLONIdFb3R/HklWMQAx3p+9w2TVQw
ngVLJPlzg1JRSZFM33hIR6zyCPDhnTYn+ySOUliNVcL8/ZoWwDQQ9DB+lyA/He+L
qJ3ixIFrLqf4CVhDvy7lGaoz6lZV8IUAsK77IiwqDiLpu13wXzpBZ6MYxzVdJNYO
biwdU6C+V7HcKtpmxenmnodZYwaEayml2avGJce1uCEvXmQ5+3msV0VgR+No/2Vj
j6srRDIQcaxCM/MNMnwigACHV7c0gidrM0N5xMp/6AkcuKrV3M1Y2rVIXOz6KqFx
WfwwqoEJ9nI8kqbWBnxVQnJTzKtutWFL2ZUQE97x/+VsxzLsxLRhkt8xhPnGKrea
LDYLgMecU392X3SGzMKJHP4Uob16KNDHCBJ/FDivkNY+VOc5Y5kC6EMJsO+0X+27
kboOnmoLnlFQ/k6miwzTrLDnHqLbEQ+/SK+Oi2zl72gO+t5KfXaXwnGtxxhS5o1j
cruCQbhaXb2YuYeZlTjeL7bxRFdxPcOs2AGk6KyjWWP791CRxyC5Vutsye/ujCUi
V7fS4QlVsbyTT0x/aynvi7ke5II7TBHlrdDMXu33ox49W8MXjvP0293lU+Iqhdqt
RzgBqmYIIkA92/u9ZeIna3FgnpakWkVyPZfBQ3WByApIGpLNKEjgdvmc35/Q7WUB
aPxaiiSHh/Kxs7t6ti6W9/luGXXn/MJK1LOBWNEt8j2S2WePWqlbY8WclvnWpHI9
O95x5uLEgHKg1JBhYAAGbe7EAYNRCt4xC83x0sHlgqTstNqWeK3f72q4fB76o6LD
Nrt4jSJCw4ffDcdzldp8hMN6/ras1DClHsgMsu6vBGVi1muPwSBcsGTmkYb/xCLf
w62aOm71Dzs5RIeuLX05/j7WtbxKm5b6kmVUQ4SCnfjfJNToSzEs0rSzrstU4vqQ
THMdsx6H3c65A2BraHUNuO4J5M9D1uJAMQ3rm/FQ1V1lxMgK71VmK+WyDsWtCjaV
F0PKvu2ZkwYS84YJ/uTKMclFr5MiPSn4ameVgLG1mtVrnMNw+zHS4P6JgGpuV+bQ
o84v+qUtNPw675klK68M++nLcwBoGFACPA6zZRWbaD3t+91NKPGNxge7ZiF7p/LX
XufvPi1hVy51K1ZYc1C3SePt6LN+jmHTXxRm681YsJjZTz6n2CF/CyM5WVvjl9bb
Ee+Q0u70IBEaltP6iQIwIWLC0xiwoj0vekFKXYvSIMIZJDXXIWQ7Hl2E9LhuHzFx
aRnuSywZjsDmNVDhpwOJHI5vXpeBtq/6RJzwFR8MpKFnKRkfLsfexahqZ7gi1AI3
lw1kUrIPSIVLG6Nwc2yIP38l1/dgS41GxiX+jV/sNW32GjQ49CsTTJmcWbk1Y8CI
CRrLuCCGZb7yXt7JjxGlwCLF7pXlup12e2p2QQilZUTKBN1yLwnP8zAbw2k5nU7D
PRv07K/0LAAsgOxI+zQL3PaiJck+xF3pDa1sF3LN7TQdK+C54MEmZ43Furu3PPLg
87X9dPueYDod0cx1mwdVux6iHqDZx7HlRtPoFnBxJK+qZaqlmhiUv5lO7tjCP138
1KUG7VmKFzO7OUnY/xq8EXhLLDaQqFez/UbfSfNDv0o3W2c3R4xSbUuvs2RG6s7+
oS6nh/12ksYQtli7EhkCz9xEQXh+uu2ds0jhJHwu+ptLnqGIJACZDVafAzi0T0m+
9/29lZwSsq3e3hMjZnX77pGQpe3GbhW/wCiYAB+fhOv7sGEp0jAjn8GKedRnwX1K
a/cESqjU/RKr9CvG5BvmURuzZyMMGVWa29UCTZaV+Y2jomalTGK/WgyxfRAhDb+D
aljlAm0U9MIg95trpRKwEotxa2/1r9AY3ty8Jn1TTtlpgA6IU9SOmwxsOKOcVdi0
MplUb3tiG/37/soRPo9XILboM5WWOycHLB1lkkSdMm3Umau0iSaurqltfnQ1Lrzt
8bBk6d5WNqAU8FDioC0vYkgEc11zUsETQW3C+vsEy6yMygR583ylHjDAERLUCgCU
kUEwiUkko7MTioOHyDc1CMveaXoLJnqYoBouq4HAmFtNJ4xpa8pjibV09pkKRM8o
MuVqEXm5NVpDqJv8/7S/R/fU2U+JXMF+3XEZ2f85CtVk9afSGbQza3Uw75l0BgHM
XJE6GnwujN3Hf5sEgeZNcTmMHT25Jh/UWvOZhx1YYWHdxgDesXBoKmXc8Cvpd+xg
maKx8mwxMzN+//yZdFgeygygV1TE2fX97yrC9M/Q96fDcIwOUI1+LnC8BYt19FUK
Tk2bwIAsjC7K2HP2Yxo6c8EJEe3hspvpUcFmvHk1xECyH+JhUeX68Af5fL1IZIc5
CvGmGiE1F6ky+HGsHJaYqdR+DwwPdGv8qYKS1O3O1G/wRhLMBgijpIx2so902lc1
mweU4/BaNpA1H8JQ6tiv2aTUhQG23+WIg4DzjFWkIlg4phKU3Cuj8YPBrMo/uCxE
bQI8x2Lz5421P3xsCzzxfTPTQ6zAL/8bobkNGbI4FFOGMHaZDtlu92cWH6FU5ljO
7imfdL3zzPVhdIBHlyhYlAsqj/TKy8OBUK3BDJH4lvBO1mEDIuXiCzK67WysHfdS
NvcjiQyF/GHCZLpmn/pPHEjgjqZwazHccXzdBCimIoNESB0SlqYPRcmeyRYDLDDt
Ah54zAdp75LAxdGNInZtMwr0wTMwOoSuWznBWWQFugFRGfjd75+G3Ifw3Wte7Zhf
hOuMTdiiov3uuh40f8O67xmPdj2LZ+MtiQemtbd05zMEL+EDaLN9ZO5O71B0Zfl0
qV0UIUfw8zvaitu6tJ0L03ZFl8xNKFANi4BpEErmJQ6Q8s/f3tx/e3G5TvU3yhi7
oCDjMSQANwW40VrBfxqheEakXx0EkIwL/RTTgZfI2PEM/KJ6jNouHyT48hovnMZU
q59t3xebt9Js8ZvbP649Xxdc07phI0AdLDufpSdYpE3LYqe/CFjPAm+AkXkfS00R
4XO4cT7PyJ96jUwlykluNfgtT2XGq7dkg5nxxVZ6yKK+DL/dylC/8kjQzu3i5b0Q
QwltDGJ0kLk7krwEyyp6JHLWfE7x4t+zgZwiorHC48aCFZ/k6eNT7dgpTdmBEFsu
9vbHN1sOrZTzlvoOLLBH+jUos9E7gohxDT/ggQJ7RDDMkLnRats27enf4XLjKIiT
aJg6uz5Km6LsYKXCTkRN1UzNcopytQYmEYsE699CTJbae9kxC6C82Gx+kpl5rfm9
KOC6GjGoVfeXS1uTy8NRIf4bNkXJkrGmhAFx5kU6hunpX4/YTI5hHoUfV07gZBVI
qm83IEotsiB5osKprAojjCj0KiUYxWezuaKhyLg6iucuJpR3pV7LTl3IqS06tOYP
TTTDeaFnwb3O78O7q09wFeK0d3R/EhhGaCeNTK8mGftz/I/+ryOeQqkvLL0oiXUR
xMyw+TbARJOtIm42HZVsWj5ngdBSGJqyE67KBJZ3FLJ5oXQrvVDFhkGi/LvloBtL
X56HxLjSFX42BU7FzRPyBRzaii6bEspxqhN9W71qphnbLYDsO9dxNCWN+xjjLeRo
p/CYiPj2aUivchwuM2PtA4r3ijJyZPxeepTtNrNF527KrCx6l+xSboxEdCnMzDcF
vgyGmxoD4xWcFsBA+mG3nXb2cNGCUFvm4C9eutIs5dreIluZu7HGwEj6Gq7tg9mf
KPwH5s0kNw3W/rT+TsI5SQpkEjVMUKP3TRw87Is/oAH3rmjn38vCJaqpZGNHGd1s
VkVeQ9IDFWZOaEBwWvjOe/SE+FVXRlrLIxaOjZF1hJu1g0H7biN8xLadIJ1p7l/1
v9yaciuquf8eo8GPbp6L+O0Bv5Z16M5IuXeIZOz63uWQva6Zkgynr5fi2xbrXSn+
IomL8Q8afu2+s20byJRJ/idPicTa1M4UwrRBnypA6DdvX2OplrGJ9+kc6s2qJ4ST
p5YZu7TSJI65OtiIznFyauBGBbAknqr1I2dEoECYP1uTBdd+RAQ59au8qKyTymRL
ebgAf8R37SXFQ7vepSZ4JQkCeyivI0JEFvtTilvMPAGg78sHTEJ1iyyMKg65+UVz
oK8fQ7Whd8/QjioiXFvi9FHsn2Vzygdm2KCtK+vZ/BQluELVFYFaB7A7+5fmzLyc
n9fxMmUfGDcYmBrTjH5np0cK3o2D+mRM7bwjjJS85+FwS9IXBzkG+mQGhomH/TrA
P1n0wtxEDk+smgtFWJe7GcFRpSq8FbEs/qMGixqk6CuMRAAAO2kMl0GbQxSMDAam
gZj3y4k/trd8aeB/JopHt/VekyOA/ByvVMvAv/xwXLLWXLi9GTm0aXZ7xSQW8lhq
K1oM/91v5fY7KhBJqcAbadVwM2T6MzFzQmR1GdaA57Z5A5y2Nwxpoazffv+OaW9R
NBzs0e7sU797OJ/1+GoLgL62Z86kd4/J54WhSL5ZvNgS0d3UfbfUTipH0yBf8/of
+IBitU0jf8JvqRlkOMsBFWALHCSzBbXqTNqVnMqugHVoiqr6oBuLPEnyxEv3PesT
eve1La57lrxinTdbkYZsZaNjLLefUQ38b+N317Zmmo7E/+oYmV3aZh2iqLW6Elwq
yU39CYweL7X8HyNOMpl9JeGmruTHY8cp75AxAMI+hINjIhLd+x+FA5ZcDGwXbBgq
aEsjpyt64P8kHJ9rgIFRcGGK50M5BzXkKQrBo5VseegvVP5GjE7gqY09tCeRqcmm
EUN9+3PhjfKFCoY5mSEBp9//M3st+7NsP2XGi/soXsssDv3sgEhB8z08Mx/89g3u
v20PtLSTSb1RFDyIXQfcmawwqt84u7enVSaULaX43wgQkPCcjRkcRXc/vFiONfV8
AV5QM9yupPwBhmUV05h/KjJkJnA8pX9xexIQwD4Gtfb0GdILVurHQK4MCvMatoRZ
h+IXzvewsEpDzxfKEtaV+eD8oAA46LGphXvy2HNDp+8hxp5b2b3wbmyiK8xk0DkT
wt2EcWnr04MsSaknA17QEvQGpPA61HhYT6XZugSIntg99fqu5RtsJyw1b41+JK8m
mmdUSkCLCBn26eklEHF0WYe/S5BNQd13KkU2kcKzXSjy+WO+gs+Jih40HCqqlO5b
Lqaczhuk6Nt8tCOOyi1c+6+4jGlvmlhKbkZvUD/2bchXCbwAtlZqPZ2W6lfVuaug
0Aq0evTAtmK7z+2+GDSsZwiERKcG9XtajC0ofDijqPb2yYN4E8sk+THoSa3K8QK7
g8obpKWHtAsJTYVa39sRUFEDh/esSNfzpq/SnFGNJWfD1VbHS1KjywXey7v9J0W6
g/GLITE0EsUkyA7AvWIDx/MwBVQFhTUAyi8oW55J8nG8E8Fd82IqBRgNhC4yJ/jd
CXzmAePbPQcD97PqzXoJbR+7RI+zW2oan44XLKXqa/NfYgQIKC22ppVMeK7gDN1q
WqzuSU5f0badI3CYSSFv82akSU0aUGXvySM2NGQLXnfUqsBFN8j2K6l4Aaq02Da/
GSgD7YUYgCH7R/+1PmBeYvqJGA/+ibV+KidTf57R1d+yI/526FrCezn8QQaEwCFa
vyabjFjub5wKDGh8nXyAg39hZfu/K63iescwE7E3EgUkjqM4CMmJ3XLxoZcEFMe7
Cu4tfLingzNcZjaytVeA11QyQXKw7jKGU+9Tqh/fkqKrXQRk0z4aS9Z+tbJRZzV2
lq6J4WHdxhTRy/sj1PNPKIZ4FKR2B8w+TK3lgTx/R+Ixkev8NZU+MTfO97JPtjpx
Cz98BttLnOVR9hxLAozYiuasiQ9gbm+vB28PCjumRUddgCMapsjBdMl/gQfbsWNA
PQqVfhPVFGrSXIRSXIVd8QDDtdvINgdWv4ibHorfcTRVBy2kwJTvqfKQTqCAStsU
iqW4Txq21aFI8E0zkT++KZeBGx7X3hDtzy2f6k11Uaw6ruBDC567plDN63JLX7Wn
J27NyZihC9TB4g6m/RT6hExCUGz/QSdWHvdwLB2BBhqP+9WUHclRHiqZ5vBabLYj
a/DI6VjTj9o78oY7FVLUtyrGRy2U1R6YAKn8iU7w+6dMbLlUe1ytYA2jMfPeH9wt
s/MLgChfXxI3ora0kefbwV+eB3ve3G5CkAnGQAZgTqmTj/AgxyX9aWOhmX0QpslD
uYSGzaTB0aDnSDQqPHe7n1OAAvGQq/TmaC5E3TnGff4lkN2MGp/249KRgO175jz1
h2bu0HmHN/byeb235awu1ERu8xtX20pQtub+9u2Rn4NXxFt5J1vGMeJrLrw1L5Uf
1euwmMAEXeWi9j8tnmuA+rfPZF3Y02Zd6jcbiV0+wIVp6ZfxJmqXRf4GMTJySl+D
qFxpUBrjIjEuhS5KG1URN+laoFY7rytg9EoJQkELK/JPTB1y5HRwGO1uLJYk7GfE
WegOmmHdK1vOvt2KMB4zam1YLJQQQu5i3ceRJG+VzXIezLs61k9NH7CH+AobqRBZ
sRWBarnh5f/NquLWqRRyEb6vkheLqxxxCakpbeXBGn0Dd4+LCTORJCaG9ibLIUoT
Y1aK/f6zd+StLl904DDv3m1tJB1i/pAV2PebQUzeJG9bEWKh0Cs9GUJz74++Xe2F
yj+2Q9oNW2YO9TMAzmymkbQjWznXeRKKZ7FzC4w97sNqYL5oOln+NH88NndPGiCL
RpjVaD6j51k/J/jfWRpphl8ad3LYyodx77iDeSVsl24srQl/EpBNDe1jOyIM4tLC
crQKhOkD5S5bOZ+rhuL9l7bauPzbWa96TPp0cTLABnFhJwrLuDncv2AvMcoTpBNo
sii/0x+Ekya+kb3zj6OF/hJHwJ6DKVFftcRenR4W0fuz9+/nAGjdi7FsJwh6Fsks
KkpeXwzQdhyndGAH5Y9KL3THev0OpZI2DbUeXXBr1gb319xn8DtIZckA0j7apRmO
VKOCsvisOQx6It4zSBSbi2PSOYKYzFhxSGD3Gb2BvEtN0IPWzDRRcsMjfSYcSYg3
GHneWAxhS9Dg2kaS6d4s6nhhuCFeWGV+9vy4klfrgA1my6kPHpSiAs6mcaj5YIGV
fTEFFuKObwCu2o8H/7EHxT65z+xorFtGZ9U+Wj5qIFSfUViI3LKYLUgkWXKJ2T8W
faxw7Q6gX0bjpKvF1y3fFpihKpQ/TiSZ5e+sl6W/gmaQyTLLx7nhpGkwGZNBKslv
17rDzLDYtjKqY/x3diTjvqYKISALaukTyWqZbxGGWhFmhXoCs0IGnosaz1JTCgPa
PMhYb/JkjFpx7n0MjS8xwrJefaUkuv5C6erJaHVS1qPfJMb8Lag85jXXy5JKMLj0
KG+uif+ehBm1FStyotpUT9ksV+WeeHULsxlmENmHk4HJz/DL+k9W5XW6sUFJCCnl
M0VA00ts0QrV0FUGPkDj6+apui2B77uGbf0MzMCOXNf/bmdkl+edmeFupk2cGfy+
57wE04mPmQET42560/Liq2yixewJyYbjhgCUMt6HP/+Vmq4qkSdvaoG4Ur7rP5ti
vB0G8ZEzywblhpbow24F3nZ8F63nG5jhlTGZItiPYMdNcgJuGuNRI5p9TNMwQwuW
ep3daIVs7JmELt2Lq+vCfyPJJTH2YOcB9HhDEOnwCjgo0pc27vTHnjAoxAiASkhV
eX97JEaE7yOULAZ+bpZHm4qMe2/JTOLChrDoBLKMyd4u3P7I8jJoQgFd/BMXbUiZ
3GrcCs3gs/YNqWXTCg5XErvLryrmY9drxen7HlhWD+EWakRzo+D6XnTGKm9WD0QG
5rfpswOhrZBfIxvt++ZLekHDDUJMKXsCcBFF8AvvVnFm0VpbYtyM1dFzt4wgdkAA
quiC//PCDyryORhXUwjkEZhuIXZVmiuK5IE49t4HOIkaR/7RGZ0fjvOfTcEqzIgL
Kw0TloSqaBFJBbxMmoW23TndWtEYNhNB7T9Xppy6MQrJKLOats+ABnkMyXf5na0y
KzUR37hpxQVlGevYSQ10m33of+G8JzUI+ONXogiOxvd98R/PlekwfeilRQMJd8V4
5zOT9xBktwS9VYPGXAdE92H0KlxZFukFYnyWhBklOJpvwoooRbQVAaj9/BtKF97E
lUztZrZFcAfRTRpohV6pDjRN6Eu77Zys43dqgvoHVMRTM9720E5vFEsJKDuce5oO
WXUTvWDcExNEWQ5yDp7tXqlYp3hMY9/bZcuQgECQ8ChI6mDpxJ0p8+aTwBJM46yR
pq3WzTyQFWOX0zj+kIChrNfdd2b8KJCtXe2DoqpD5QcnPk6C0p5B4xdfOl381BTq
Y/9Ilh5UusVDDldthehL6CIZ/H9pHWawqtYH251G7c0sWau1dQeflvYMiOos5vLv
l/lqUHO5iLGQVy8pNFviwVI1e4KbRXM84pNoTx2+FvGgAIo5iyHsRTGYwJyu2fzY
/yTKOhUThpBpwbjooFxmttVng7kXsl7KeVQpTR+ZDEfjmEUclxUutL1IiReVxhJP
qt/bW/b2mV0MfEeELWOI06MecmIf8+40AQM0nDmvyRxK40pKtwKtKIxqM5G4DjxF
mMMDPjqiJr7XQkKJuWbBQbKFnapHOMF+A6w65sPwzJIATNsZkaUaOinBKEkaXZms
BjUSXMm6kxPlDpsUPO5SimK3MVTGTya43JNydxGjHLAVSGQqK2424lctXxAM1/2a
BQeYE8w9j7C/rRIxfVR9iChNIC+RiH1DOWrAY2BLIRvd26jc117ZNW2N8iXDfPSQ
I5n973t7/QK5zpuDiqGl08uSisoHpIQBZiBGyBtf23ILo2emcVD0dS8OVMYC6ex9
TqotAOcb2cYUTnC+bxrDAL4qlM8TEYHZYFNcYnOvj/LoaET0OPYAOPQt7UiNY+hX
GHFkZ22NCyVJS+mle4VVmkIvhu286vgq9vgw8t8EeCWcbq75Dtw9gGBtIAL8xqHX
TdF5BKe+/oMMqBj9Eax3YukbRslTX1ol2xTCVF9xkIG/cwTIu549V7+39PReRVXS
NPcmZnizSwGUqnjgN7RWstwmH1fAIsZ4wnWvGDtycTHrBHQ8sIm31kVmddLNMqLC
0Rt5cujgZjIQyfCPNq4LQ/w6Xa1Fb9q/zfcbWnEs9ROT0juiJwJTAV9ciTKuRXL1
X4sBm+VEBzIMGTHVpf29lfQTPPuPz2pUzBHOqm91Qdw49gUPYv50GLJ1PMdObLAM
FeA0zjs4iZgtEek0b68Dugv3cArRF34u62Q+RDyKOXBuPTYXZ8abNV8NV8A1JDoB
jTz0zGxoH2aLpUiccPVZRm9BFpc2sKsOGTKTxjFEsPGkYeG4U10yg+v61tx26tR8
fkNDYBQBj3LgvZVVdEk5sKFCPuZAr3X7UHhac553iJcB3cQo+qFpXLzqiPWcD2xp
D1liMZXvSNdQsgNhYng0XdLwFx2SpZJ46vqbm/4iEZaoyNKXIJ76p2ALnI8UXCjP
5VSNE+7KKSAx3ZavN/hJ46FjJWG5ijfp20dff3TJkmb4bOkTFrRuiYrM9dqsUy3F
/Zg3csw+Bo/Oqr8Dagc7hLwVfUOI31dWXUyN010jcElenqdfl27O5yJfL2c9u88Z
bDJ1OYIx8lRdYVLizY5PnWO9Y4b4KHnikTwQ06p7H3lWHhiE6cilyCBUb1X9NkL3
b7kFLpqsYvO9tRjOwslpJSKhQnU1Km2Vxb6+DftyqVYCu+x0LAK9SXXVouu8aDi9
iHfLurdXV36qkhzbOitpdkNryewBlk4tsNsKL3ulHA2U/g4QSqwPmroZcuI36qEw
GFdekRzgNvx0aBQJQRSnbftkueBnuRJ035UJjfRyBJqE22sand1/NKN5XpWMcXjd
4DF5rSuv72HaPt3jFO2WJmCx7e41TYXmNccc+G8W8Uaog5mnYUmhA/An+so8csUT
40OXlLGV9WbZk3tmLRq7dLgdPpmPNUByEBS26flZR/oRqXS5fX02xDNbns4tpmIf
yNRITjQPvYrAFVqnIf/T0i+78PWAshax2Q0aBGfVdxTtedG3YjX0NNDEip74qKY9
S43so/4l0epEvvK9cZjHApSEgyqx13KKqb3Bl/TIzlfgscqxkR3HAWwse+mAf8GU
4hdELkt7PjqfP0XkdiFz69dA1/k3tAl6oLyUMLFQxawkg8Ufcrj3chN3e9IDyCSH
u+g34e/32kTRxW30r6lmM3pbR3t+Www9IrqczX5eMnC1fMEfRkVyGl+34lQrjdPz
Hq85M5doFMSetdBlEvb+tq33lEo9wyJVQPteP1ZL1WLEc9GAUuhkvgEwDJzfycIr
UVVVZwd9OqUy4FzF5fGNumw/+uJf7pIhbvdDBNxbqeOlSE9MlgOmBebWnjBUYJyN
xrqFqMFy61cCcP2S0708KaIdTAexc04d1gGUZrrX2S1VyvbvQr8oY3nGInarVscO
xMy+ZgpN0tWVZKRZyV2jK/Iu1fjSQazTH0OvTZ2CCYnEFSV9f8tjo6ANusxXJsQ6
fiJUvSWKhMT0J0VPX6dyfn4duLU/VIjn+GUNK1G/MTPHM6etXoMaaHKbOmcpCHLG
hZfjrX2d2gucljqZtjFnjaiBHHhJnu9y6nd5kek+7VbNv38PBVrNCWHkSTcbha6d
vJrCSv7UgrdDfMJzm82B+SRyKreqdnlkoCnFaY11oHsAc7xxRDQ+qp52a4ZLQ+Lc
90KEx0Pa2e9Px53aK6Z+uvoNSUpOS7kMNIDYeB3CpNonzl7/htArJ5LPImjBSnyH
fS6ZEs0QuYGFWY5dc7OSAMDGUjmCQxJbks7OFclPmWd980Tk2JWiNrsmDHj2hH/U
jp4hjrhwbtfTH1PIVw1Da6q+0ZCvOnrkvy7Ntndb7znrgZ2AwBzCTmP6gQyljlgn
jyWCe3DojRvt47X4JU9nBpcCb5zXI/551AYMvBLZ/+RaObl0wMcthd+s7cj80Zbq
n5XUZ2UqwqJjRwRQHVmWjLY/DYeLLjgYSvfz25bvCSyqDkZN0wWLJyKm8bXcfrvD
JUCsZ8r+Qy9HlIiAd+ZxLLvM/fP8rL8O6FaT+XdJudDP4Uj91wOlDoKokh+YT/rO
B8injLEfQgCdXFFdZSKFtv/TGlL755ikqcYC65vU5KMqTp+A8wj5ktKfZg/G3zZk
0CkOozFr5lnDTV1Rf267A0Q6VzDi9+tGaiGf5ivnjHGUC3xZAscnJpLxJ6G4lDOh
GQttlk9cwQn4vVMmm8bJdudX3Qp90urH1KjTZT4o8lB0cSuwXLwGd/nqIMuyVmOS
jz8vRtzDWY3MIO4hknZpM0miUo9HQiTGYwkLBYCCBGcl1EDomj1U7xeZeDhUrazv
E9FTj+yla6WQs0SSsRwm9l1gJRVbe3BySVnAGq/QNEZkW2fs8iTbOsYa6wLOElLd
GHgMLjeW3qYbdt4WGSVR9+9O193W4rRqe1jD1U0ekAsZr9tz0VXdVPqwFmgHfCGs
0gK0D+EoHfLZz/wgkSATVt/GBVSd0UoZXcyHoq9iwtGUx0QTh3TmV7rDxWgImWf0
aeDYYKWHbZXI2h+/DHqgMgApu6gv62Kn/C5keDM2bdate/7j4BRE0lmV3IpHotIo
OSlF2pMrXQ9H0mMyp2AWnKjYAlpnQsMrb77AySkOi7GOFwUho4sZH3sgatqzgcVK
y4oI2J4kUljczcHhKnpX0I6pdzytjiOzOf+5gLjQ14D60nWZzEK92i9P7UtAyDl2
nVNv69SNNV9Uyz9wgwk5uwgqmsSk/gEbB00b6OlSpj5HMGdHOWrTm3GyP5hDkRFJ
KiOfDEapSTyDcANbEo9+fLetxRAdBMrOZCsf0N5vp5SMfiebymtLhZtYhSJ2iq5r
IlAwqVFRwYqda7PXhns7gEVG6GqK2JPs8kDZHIvN2gmAM0NCCerbwT1ebNBlZ5wU
vBYdmZ3RoPFSjdo00lOu9gJ6iwN0lMUKEbRjbx+YC3v67TuSiVCLyQd9Xf+d/FgG
8Xmg8MRsCGO4feoUhmOipbIkTLsGUShGUFrB0ehfdOPpIuK5y6U+5w/Jvp6QZKvv
SfvQvv7hMAJZ+j1YMJDpL9kEebblWRc1gczILMY/hVUhocmaUYPajd6u466glG3j
hryc/QAbDIwathgPhfPf2TrKzeMBtc1JQI7ZNCdgIgSfZ9cr2bWTDEjAHUn/viad
UcdrC7lL2Elbo6r8WTMVNmITr60D2tG4pnGUPz/g+3qlrkM7M1LhqnwuKsh0VG7h
AjfuuM2EwqQ6Snd1VvfdZCrPmpjlBDhwuV6nGdAS/CJhigtUnEYqrRfCEY3fcjD5
frtlArkPsJzq2km8LMcDXAUn1912EwGzzv8u/8+vedBfxcDKKE2sZgNLt6NANa0d
ymqfNI+4u2f7Qd16dPpI+avASMM1J93HsLs7kvxTxSoK+2znYi9s7K8DhCeGt4WI
hNMl/xeQ/ZXm8X0tu18KwFujCn0zksrW4Hm6wS3JwYWCpuZFxhIKBJ1o0YPKNZFx
cXrvfRbvsIQ1ltYuyEDeuPyoNRXUHGh9uyZolAIJhd6OyZ3VWSvjQN/t35XgFOWP
WFQ/bPKSUmqx4/w9OaKqRxKxn2Ca4rjrmiM0wnu0XAVKEHjSGwXy/9v3B3mkOnbT
9h2Gizoye89TNm3B8gGG+XP3/U0OJ1f427CxQ2yUaVqR3Y6wUmpCtEEn/J5YsmzY
eaCmmWw4wKHPTefRNvtxdg8246WyIXB3zkaJYNbpfkefrfuPpDkz6lg9DM3Bpb/0
24SdL1n769/M0K5+HyOmHWrrqTlhRyPXshtEAh+ZfnBDuYpxsfvnncfhUxiaG2PT
nNOafYQur6v+fVOGGrEopeRv7LV4xU+YF8pYBFZAiBRYN8YYLk7BYDjiZA00kvXC
7XKWiZvRcAuZVddAi9xc8VIPRqfuG3QyIpqMVzqu+y2slaYfqNPg1z5Zvb0uGsNF
C7HLkwxI0H3iKdo+SWw+eTZhLicIhrr83ZjlSQJ6+GkX67gGeJkzvz1BnwLnnunc
6Kk58uVISU1vuRmnlmyrcrVNkP08vD4Da2fzSat4hWsDgUrlwCcmoo7GCqXprdiK
p3i3lQTx/PIPEYJtPxxklz27qyddLL65qJJedf3Psv7HwA7hS3orzaypr9Mr5/8J
cdqA/pyUdIKssLydxh+tANcCoDkhPrnA5bk8tjq2PBDfruuhz5Uxy9C3y/cXB2/X
DgevZnGVPfiUjnLrA3PC3je0xdZlEqX9zMRe8ciBMfpdaOJTyEzzyklBBMZUiviM
TrVBt4LW2Doa2r64xxl7B554Pj1ZRO/HL8dFKkQJbEOlGw32RdRsyKQUdvYVuAnb
2ob8Fjp7bzZfTWyO7YqYAGibxim1mkz/sCzFbLobfV1kL4O0YmVFANDHIgcN0mye
AWHDBzh2I39cf9ufoC9zybNf1Yqs2EtbhiYGcEiVAzxK4JmenzoJNMG8JTe26JZy
zUzl1NZ0+wW30lIt/i32riWFMKUy7mIcHUrYD7MVVe0FhWRowFj3pdCf2znaYb1d
+bj08L5b+3mc0M1FovjqbewbfpW4brIQ6Gkp1mZ6hepkuoG1wRIxVomdfxLfvXj/
Zei2LlUA1Gp2pbfh/8I6cxu74Q1tvQ8ZyuVWFxVAFgY//TBzF5tHvzfyo07QRN97
vyF0GW8+3ImdL4HwdLidkefJAIxJjf7eKcYBigwJGtbQR9GXRF4YB6nFuJRGZCj7
tFpFcaaS7NRXvtxExgRxPX/GMnu+SUYVhGbPAVLdOVtxNFihO6I/S/jt5b/hSx9b
fIWSmYeV8P3uBmaFhsoCwGDKVpZPn3IuPjJHytj/KqYTTn1c6wXxZS9OVdaodZSk
bEyGMdrgWLzBchRSWTmBnAKoA9HEEAQ4g3ViV5tDMGTIjWFwtSdrID8Tq554Lwac
iFbcpbP/Cvr+ZoG4Yn9z7Ld5j8x1T6gY1ZdS26ppA3ppUntpQKq9FMzwa2XWCfb4
li5AY70TF5onKJ4wmeI9VgCAjKoURuAfTxLANhexXvGbRvTymWPb4fEH0hVhaOL2
4cIhqMFx4YASfwFZfw3IAxv4ZNvoQMXVMTvrc3KiUAPVTxaW3GkLwR/YVLR+ZExL
dd8QRl8MiZXDIkL1ogE9QGoOmMwBMUyvVMYgqUc1eRjM+QiYI7PNxjPgY1CHMcak
ZH6mH/8mi/ErHzt3ulwE7z3eo8hGSbhONGSzKZX3ysmAyDiJ8+Xe7bd6mcbRntCN
9YGUCq3v4t8q6TMyt7wJ7hf8B9iu7F8oAJSp0wDrwnc8K5zSn9W1vCMRMhSo48Fs
xJB2GOUHbMDoaqGcW2ypHLBwK4tCx+1oVvvTAZjf7fgaBcg7rTLsSFlh4WVe3kh5
uwarZj9z12ontiT/qs8z1zIa/EIkUYlUl3s91JowHiklkbHfg4YOeWdxKyGFkfCP
wC+Bmbhni2E1u17ap4nUywSTf7wiJPhIqenv7sZmn61kCW0yrewYPv+Mi1/nyNrd
Dyw6iOF7t8gASa79pXKmi5EBxQ8NeTdiDaBJYJxu9ata3yeXF28lDA/ctdQcbm5r
Lk6EnzyjjmtKO76KJLAO1oifff1RsVUV1T0AUsrzYpteAw7pWj0cFWxO99YGc13W
LfLY4dYX3VBnmtTJRuNk1T5Mzzg2f1V9rjXcdbDd9iLtV7IyW+Z4/olu4F8lwK5i
geXYf6Pa6Zm0/0ulRGyKPW6YHfkX7K1H1Ptxp1xb0Z3BotduIwPvwPlP3IFPQHg/
+KJrbXninrCjprW4HwcototGAifkrr9BO7xsqO0KxWg7vQRXchxM/hxTA047E24h
FdjaNgcEQoW0vgn2V/SkPYg+w57IAujop20NxSBnyQfwT/UE/66pbZEryqzuccm+
1xQp61Lyr3OpKXGbTduL5YvO0ZrTHA9DWanjecgLSvGk7iCQDAKruJNUdY3qBpN4
zPcV1Z7bU9e1woNZh9qzgc4JUBlsHk8RkhqDdz92WEhS5LBKj60cDQKKFWaDvI5n
aN00kbsoZWdPZZh2fPCZnwrem3O0PyY7U5VlHBpBG60owcDyNnkJ79cth8GOruXG
DFqISbsiJgDARtbwDxluUs+h38BY6D8c6DG/Y5d18EoEbJJMeQPpWuVSwJvfX6mh
ZcQcTzIABRwpyPwEg05Q+z8FqnaElO/w9eqE1ejJMXKexIkUggeN68xI0nP0qT+4
c78fjS0YmoKYVVyWVyEabEl1ymA/rBI1PKgkTR2h3k89Eugkwts1rRMAlQ0zX5UC
HGaR56EJsmx2oY3XecC+rfS9HHMkWSdB8K+cgnbhan+IRNnqrdraEfqQMVTgiyF/
WT1JY706Pb6wYxHn27uSZrDgQWQ6KG8K3swqZAimAUXq/8aJtcxME19reCkRvHR9
arc+gDMx7XIBQQHIRtnHgLx4ZR3FfnddHbnlXJp7PrUtuP+bfkEWvU9jupuqtd55
xIpzERc8nsI8f+23sruMj4prtlG4Ikps1OzVXvutiY8sttpSnjdca5hbaXONuZS+
zaXE4ooRQ8wCfYFLwR/bjSJesvxOxhgdRKr+XVZ0rmNRBOTh4MWP5xWwfxgU8U9p
CSpvjH4Ua9iQ/cIZ892S5Znnv3eXWG+lO+ramB1TCCzD+CXAkBl904BdfVtXJpuG
YOyr2WaL1r+TGiRmxijRT5GJ1zaggGTiwnh8Jt5L7Odkq4wI17YKqhRadx1nbG0o
nUtbovNtgF40tpTlCjmGezvqLRXdldy1w5WzboPM8pYefSq+nhwQ1cP5MiSaxg+y
4oEPwsOx+C0N7PH90G1Q+azjW01yQyDA0YBQeRb8gvoHvEm04PsUfomc/lADW5yf
YbO7ABR/gICrO4LcrIuV6m/i4rIwj1kOkKt640+brVqiFfMGqOACYKdn5/HbhoiV
bkw2uEhTfyL3Uf8gUVc69oAE60SglUERrWbSA7zewwNNgg0DXiLIDCj8Ba/LqVWJ
zNNeoxHXh0+akKWGpj6PRP0V0tQptNDLLwU2/Lbjq1L+nkl8mtXI4IYvnkhfmCO+
+znWRo6xWTAG2fmKafPgYdKQ9iJJbbH/EOLsOflEL+BqAkaB1d1eujQlYQmaEihE
SWzeuItDwagKyo/GKNWIzk0KWU+UQxxbd4sLFnooFUU8AldVl8aGWvTX5f1K1Wb9
w3MLnDh0Rmi6hVawvLHOyYkaAb2b/Ut5wNvim4ZyXEDXP9e+YQzeebrPLpuUQ25p
Fy+xWlkRswULXv1VJzcgo9ifNu/dJnsf7sgXDFdpViPWIfQ/AePLAhqQpLNYIwhe
yFqFJkMhsu3EepB88WW/Gj42tfmkNF3GOEK2KHeGEowsl27C66MMxBPUAliC8hfk
k9AZXQMtg/GaVYzMgkQ4EBTHvf9Md6oy2nPcSn+a4TxNmlmSKxUa+GxdqHAmRR7v
Z3p6GPRyYsIll/VYP3HVcaonuyeRyc1mgOCFUymrxaBrtj2Gx+RQCF8jqyQ32Yqj
Xw0P6p6eq3P54oD4uOjywIWByFDJ5svooHB7vKlL1q8ZFYSDxVPvbFOSUkuCCbSo
yZEit6icuqG7CEUWlq/wzUQ1/0lxI5bwZe3skyvIksA3IWdn2sGlB/s1LOqhJ9Zr
1p1ux5cD195nxc+zvwTrquNBWycWHUYWwL8zOMiSk3vr22O+LZ6IMOwbkwtj4MG2
FyHlEpUmgQuHtSCPRT2EXgitHn6lmKRYHbPieRdISaalf6mqyG1NMeEAqem6Uyi+
Qz9d6vLo/SCuBov9OOiUzSQdW+fBiBhgvUUktWiWepl5FHUonAvEOSQLwMKOr5Nt
OmcU2EEhBtPWhCPuH26Io6qlXd7SzoPJmfHKpxGxppHwtFnFAKGMb26U4u0kZTgE
lU52fA9WGB5hDMWwdGrU+RRqpdfMuaO3zTE5qFHGfYZu5PJE4T1ss0Fa36shaNzT
YlojpXov2k1m4yvPmBZTxCnhW4mVgp7PIqPReAQz7Zq/RK2mzL13C62+G4yes39K
0jnX494p0FnB3bSBt+8eK5DL6bLGI9kDi6DYFpxPTkhcL1Badydu6DAbWxKm4B3A
bZi8OisM+hpbiOmR/WIP+MZreTGrJm7D2c9VSyGQLG5TlPBuhrX+Zty3lwe9y28E
wk5gP5J4DQkjS+VrxO1stRE6Wezlx+J9JhZ9/+x1twQxMWSRyDYsauLNtU++UQcM
WyCFDJvuXQ8acPXqEiIn1e6/F2xe3lNFdpR2HFm8HIFhNVEqo3ctvZNppb3QZiI+
Oub+xE/8SXk52ZJE98Ux6+bscz4iYr3Zc7rGsLvPo/lN/IQ/sM0ujjI5poRXOWur
zPsWHYJXUnrUb2tlfmvkFzvYbg16Ehm2M1fgjuQrdmZvHz0WdFovlSUAY3uacf/k
Mwf9ioBKa+7PmoW9372usVgglq3RTZ5jHf2TOtPQA2DtC1wwBvaHI81vKIxxEOiM
0zBPWNitPnCJjZsElTZRbfrEnZb0INO1ziqLdUQBxbpt5PMMX/fCh61PcYA1avtY
mG6LCzgBefFmbyWhCxC9b3nv2+/Y/qwqY6g8M84+ug7aRDT4FeFQu4nJtj/ZL8/D
CBMK4b7MlZB5CmfdLJcTvUOeqY1kRcwhOuYBtp8+YTjcPH3T8bhuzpS2BZvnjMZL
VdkslLSHMn85cEFoPhnP1fblmZSYcqS1sqnec+aguldBF3PacJ+yyv1+nTqxCJFC
uHQon3e2q5zqVoXvgGAuck5dpygwH/t4ovn0pCkupmUMay082wsr6KrjFul/JkIO
7I704CW/mIJlDtD7hAKzxlhryxWmDfoIpgFK0lh/XS4KEy7D/ZBmpZiWF8V/y3ol
PynQ48XDrhc1ZwyvnxhxDKO1AV87wgMuDOkTGPabB/NeE2CNtidkEt2qf5X2Th3t
2hlAWG0Au04bKTOAbrlGB5j9Wkgjl/z+/ZqD3Ge9RTwhwBLQJuhWCseawl2G5EoY
qxfdtAHIhkIIby4ZgFwev7I0n9jSuLB1VHyIjynjjFnbQ/gs2FfkWDvzSHUszrT6
uYKvb+Ab2AdyfCGNy3QcRwghaQvRKv9ruVRWbTAuXWIgYV4iWQtpK1yZ8iOd92ss
jzMiChY8iITT3viRZS3kSKlT8Z9pxceWnoZZkk0AQDWLZQlQTDxaH/kOXeO9F90F
4Xqng7JkA++MOZy04ped8HtWDS/7b8URDyATUlPVT8s0z+xvw3el39MZCxYn2bUw
ImegW2i93fkEDAF86/dI2bwjfheQ7BJL+0NghmFzZ4XZS/T8bFkc0ptVHrIo/xdM
IEOntIMj8HE5AH8XM25jR+p4xgbzUqp/t5H7rl/p/tFx1LI9HkbhDNAWDh2zeAqT
qROgXmBuxiGKs8zAvWSAVVvBnDJvTKuaNN/v4Sz7fVDNwD5Cr1q5br4ndhBSooDc
giYTtNtMItBRvPM3DBlSdExsbs1Gl4TwE74mNeWbfe37nqYdwB0WmraiblKNV/Wj
0B4+ypqI+zCg+y9TV4PEVUCd9APLK6h7IvjWONbJlGwBMpBo5Ac55DWpEVlN5wMz
MeTV0SKBFCOryxfjPDegDkV/YPc/LOJIaGXeCgbuYcbZAfnMH+0P0thISJruTapR
KtDGJB/POMMAzmNQv7Za7NOtVLuwpBrqvnMhD+QzoOD0RXzLCAxWquVyPFW1SegO
qBMlsm9OGy/jeTuxACaIauu1TkCckugV8ialt8QAC73zaDRpgL7PuC7fVt5RfxaE
ADjjUA2VyrHJmnfcAHNQuOLGsHqtsZuyiOHYG+wgLLBIQjfEksYy/o8Wp9rsZ4vW
jEQL9o/z3Qg9XB2aLab/uCAKST2P/ADJEadUAyBXRqzG0oKQ9ZX3fLRZUKHnhhCW
dxPN/OV4nbeqdpwlVi8JPy/p6iBW3z06U2+EXcuawoIECJu0eGrCMDwlr6gB6LsH
lY8MUIWkPamFJcvOXFssEL5NALc5TUcHhIi7X1EWTkMJDhTIVMijbqTjmKFTDKoQ
P4PnE2n9D49J6PeY1HmUv69XQ7YIMz15uLGjCpHkD9XsimPDsntTTcJaNwwq8hfA
UeiTJq9LW7mp5nRi+b2lR7plKmSIHITP/auUKJYnzhVNd3g9YgAvLeKQ7w3voEK9
anoCFwfQloHpAOjesyULVKCTirAre6gAQDn96M/DzMYT2h2gGnJ+vVAIa2VVP28+
Iy7pZqi+TbIp2CiBhwlH8VyK7HKy3pzpT8H0T0tG8tIEhVexifto8yHN2PniOfvC
FowDtPjdAXYmrFPtBakkv9DfMOaa9AoMFUfn0nbocxEj4vqacomqVY4t/IBNCuyl
ft1sJzn4ts2/MGDJbe1sIyf1C0NEQO2CqF3EjOlv2ykhW8EJWaUkcrVVDsPuL/99
PxgBc21678NN5O7AXcnIiiYitOeb/B4VLKd8ccdsrLSnLDAkK3PGb49y2pR6llrg
5KqpbiAYEXkYLhPtgu9Rztarnm/Ddm+ZiSqVg3zjbKpdkWXy2HtOCi/87JSY7G+4
3GJhkO7BpFjdPWt91zctYT0q/5/TGYk71Nlr2TSZv31P90wcjTCdLeyel6W5wKSI
mQWdMihaGH/5GjEtAJv5BumKox7pW/AqQeWrc9pxil9jarZVbhTy+sRBrmdc8Qak
pNPVsAmuUq8dZqBSZNRzIDhFbohyv4/G8rBCqMooQy4x+SfCT6dk1LDvxLC3+zKG
8exv5dTjSj5h6IPS+6PPvbx0c3HHppn31Hh0odAzKGzt95w6UDFbfyjtiH4bLANC
7hoAZ/66TZrBhOEEqlBTv+q5PEqFoRrb/M4qg1P6DMxc6OOQuUdpBu1f7XHJeO+j
4HtKVXhpK2T4vPRJzBui0XkAj2fpnKGn73ogZivAmpKfoqV3TUbwWo03C35rWxQ8
+8xVTvqzJ6x+DWi3tj4r65XxJlHHyHVXnBabZdlK4690CCCQlgrggyk4SNmjxccD
7hzhOEmweYXinkX1XVSZjRVl70IBUSAz1hiOfd9faV4OFtVOOfIkD3QuUk8cWw/2
zOLXCe9o75fWjnb5ESkfH7lZyx9R7NAsQfLU1vwZ+3jafbbFQBlk29DXx38CMnTx
0aOQkeqkxEdUY+WQ/T/0Z8Z8u/dhJu0nH3Kp+SNSjy6KBT4n4UZvGRH3P3/i/P2G
xWk1BXbHKJXa0bCpGn5Ozy4WuheGJRD28fZz/6U3DhHaprTWJrjmfT7NC4Pt6nrQ
6XHzwELTk4meoLxuEq/yLdJkEmBjqAuDge1g9S9Jy3cjTAh5mzNR6hA+6FhYe4Q4
hzICLDUr5Ug//DRau3WHNNmVT2XkWPFa9YN0j64mDHHJvF3r6T3d8CC+PuYUBBjo
c8lPMbnkI/5j5fiMKOdZMcKYCiqQtEVs/jyy0TJfI66RrSde4gkT63cH451WixRV
+/LYF1Z5PIMXGwWlfV4byPlnNmPK4whLz3SBB8E7YFw+D0UnQZdgG71m/Q+4WLje
TBHGHBdNWb4BNQIT5Z/orUE4fmjOtSp+DuFPGDch7bDOO9/24I0PPrWqyDiHP+BE
/qtrIsP6ZXYNIPSQOJdb4SWPGSsi+vm3V+nd+7YCfdrBVEmLoqDAenYMDqzGXY1z
a5G/Q2o0lLFhcR9hOoBVlUFHFcLuO1i973q1kXJHBCYZCgFWlBCPYE7ko8hMrewE
asu6fSx+FNifpKpptT7O6n9XL2nT6NrVEzbiKpExv7hy09muNyMc3b+Os8ruXUrA
nFieQih73e+qPhqHVHtlWB7+CybZ9rZPd2/nYqh6Pg7J2XdTAZsYeAabpp9EYZp0
NP5fUl2qGUTVE9DcAfV/nrnN3LvFQkyfwZz6rdcwyVl2ApGBaZj1yjEVsGEp2rem
QW7m+fjiShhC9lxZRjqqxWZp0W7RgXL2AjxX4dz9SKoseXt1ePq2RYjDtR8tcvgs
Q1Gct1Yd5LaqdhJgTx6DhMgdekGwVPDfuifnqz3NixfQbNP/CHFaphy2R0yRYnir
I7wB5sA01hrHBlAHvQC8Enu9RH4nGN87lklofeMLEBLfaFTdz71Kx9orrT4ajBo+
P5ICZWTevmbR3xuIwDUjLksH2cOyMO8IiA31Kp6k72ZapxsTEZ7uEvs2hq09Rglh
zkcYJjptldKxpwoqIdgFwzHOWnkFRkduvLswDrt6luFRlEI+0k74MudqD6hMWPWD
DV2SVNgpduiIeVVLgao9+ePjGvKYv2r2zGINmO/tDxXi4lgoT8an5gGPeWDEuBFz
eVJHmJhODzoUXKerk3f2xmOGgCo8C4hTKC3Hv8X+3HyONB+MJw+BuGa1tJaFStw0
E0eM88wjBtfk6P41+MnCw7HOG4qqiSE39N1402hgbmO0V4BK4CphK+BHRVJgSmAQ
MclRfVv1BqsHQk6B7Y7wubqmCTeR5bTnICI3HIpw5kr3kGB83CEyH//UkQ2FJFkW
WMAG7aWCBLQ7YWkSm9oQaLw6oi+eA+DlfgW9A+1VyspLE6K+JOSLzea4woiki8E9
2X4lG2WsJqZdiPc1+oWpFf2fv5lgA5Da7IGHZ52OS4r90OSqvi5yDJrKzyo8M0FK
JOBI2w2LWAjYk9Oak/yivCJEPEOecG650KFzZdJcw4FbVZ3So1iYErGhSy5U4TrE
gD6LI3CzLDFwxM9phIRYbaHLWiUbscn125Z6lgw7h1yjna2+Zd8Y/uBGklz59WrY
HzE9GX/qB9f8O+eTsdVNkPakECEuwc2s9uCIJLNVdK6Jnf+eQxN9Lo2BDOlPk+pA
nGgrw4SKkcjZLtPnoRGMNKXTb6/7BnMmM1Ae/hmQ3Cb1FuOzUNtf3AK+0s8qvv+C
WIGMH37QirDuaPJ4PWULdNWTb4TWK+d+PLWkt/cBsAOidy3nYfeYqSML8vajtc8/
7l46IIi9kVA4LZBAmCGek4SzfLfH3ictBgVdSsmVr00brfWAaBjHmn/LOCCYzu2N
lH/p6CvYD6vcmTFYgqVVr0xNFNarPakSNXuvcYgiN0bV3IY2HWwz9VxBEXP2jyUd
zXrPfIHI2HGcLrRrm0oM1NFRQRCJEAHw2WXqES0Khrg9iBi1K8lP0qNQEA5unRSl
DU8ALbpgSfY0tloKhM/CjRD6TssxdYWzA51hQzYDoT7OXQfPOVagUdm8pNHnGD51
qR9P7IhleiV0okljOI9+3WDEa8T04Z3dxvgxMt4rxZDqMYpcWMSAJ5uj+QbPPqoh
iYwkhKLxAaHUpTqNqEbRjPrYIg377lpPSyfAYV5hXYF7n75LgVDBWhnPgIYDcxmz
ySJDxnYgJsKKgSZfVT61AZ0uZseVgMuWP4E2GO3BrSmjRS1M6qomAvQdNqX3Yimg
xMkEpWmo/0MjovuaypAKYjcAyd8toH7De4XYMJR7EYN6O3wmNI60JVNLrixjzA7o
Vs+CRS2CrMEgohqpu9mpuCWO1o9z3xohtVpwcqzOxRmV/uUB8udy8hsYVo8/tr8q
/diRIO9MIbZX6OvTJGVgf19LPIy7MvrkkF/oy6GYczftorw2nXL8/oz9J+sw5XuD
FQLWoR+kb9Q0F3N7hqkHKgkOLnQ71HH8UoP5APtunPZ+8n1nktY0n6k9tCn45+ux
hDOn9YGyiWiCSXnX+mhqtjA5WYtACyWCd2yy7vjDZVq5Q1hQBHzqhsFW0lox4H80
b7uViy4NNfh3AjICUzzuBSgbp8t6ZoQM7uv6OFMIY3BtcBBCLCPSn/kcls2TKE81
+mfJBvatqIX29+7qZGttNUfliN9f9CEDu07nm1WME0231zSwT2zet/fBjlb8nHDA
THd/ZYHc3YJHi4vwmwn6tQG/UyNepGcOsxUefFqC+ySoifW6k8MZoyvVK2eXeInd
gm3oqYT3bAkT27W3WZ4ChbsTpbfSfCicbxMFavGKozQS06f135vCEhoBW7fudcqr
aAhYc+LYpKtXPeV0IpFxPD/ZW1X1sr2JxUpa1O1r+q2QLfoGEXs2diPqkQhIdu9l
d8a2dpN4wNz5gGr2Brjbn1sQByzCSxXt70g+0OPzyoDutT9b2zMyQFooKuybZ3RD
6RF+7GGYuMFqr7sqJjuaIk8ue/x4/qJKccM/l3PGAZ9nz4URsd2ketKhsCx3d2V4
Qgm1Qnp2aUgSUXb8bgKDxF0iNsdjPcsd3UFdiZMbKSjOP4jnFF4T3rMn6UnsDLhy
vD3sSG3ohd3Z4jswPEZvm4nxfmSnQ6xgqZVBS83H9Dddbyz/mjnf+5TE9Jn1FKP5
fWS/HhJ0mhHH1oQmW2W6aAJHusx2FhF79Zksj/jYpwNFhuNY0dsbhc6c2jfOSfiV
uCoiU8w+STgWCktuz2grBxmV+rjUmZB/B7KEajZzROnTCfiLpKIqp5Kp9qQrnviy
eTFXJ/bql9AbWrbCQY96kW8/TAEb1KnkSnlCBUjFBPWTElhAHPSI6VJ/9c7pveZy
ii+UnrAb/om1MRKP2YX1uls2LouFcEEJkMQfi0dUVxoEIlDmGnJv3JT1o8e+SBga
9nVQBkOBn+gJy32R9xAW07CrGCRYQP4GHA4lJ+Su31uKKoTwncJ+hmH2js8Ta2gy
VCtD+pz4PpwcMvK/QUt58j3L4mvX98ks5AtdJs5HQEseVKvhTxlZPXEKK3y3vPSc
YxeSDoYt6y2Pgt8a+kqJFwhE3LdT3tY1SoBWtHyBjz79KES4pJlDrzJINXtjDLqz
4W4Qi5t9i6AmawOKqeecK9VmReNdcNnN87nc389D8GehGmR4lgCaxNaUs823I0bI
TqnDKKiZyQiVe9S5ijqlsBRu1Ddchnb/Yt60mInPjbliHImrW29TSLxnCH6i5bDG
Qoj9PfAkXqQtqhBj7gY1aboQ+HLyxuAw8wHW9+pSl37qegJrBqpCSrJeGjc5k2FN
gdfcUNWumwDdTSJFDaZiT1b/iRfdoW79khHjV9QDzDVtlN0ZuQvfFXxWZafn5oXD
kI1JtcGm68BWo90DbKz4uOEjtryE9dVlMOGf0mdKysQdwOaYLcEv7iIYnsG/0bXa
i8z7loNZaD1SwfNSqpx3SnZIR+pTsErzpmtIupRtVrksXXetMQGATcXJoQFyjHDU
kFeZTb3u5mga1kEu7bi4G2Jai1uJQaLflayWXet1pRRVKQJkwjXxlIOQIOd5UMIK
GQbStdkBn7pu1BfdQNEfaoq6Y/l7E7Eu3FCnRs/kYK2ER4YQJ+Z/gcTi02oSekJ2
PfjEXEI4uz99U/s8E6LjtIW5Ra4kY62qpDe8m5BGzVF4OjVb3six7I/SbMGQucsQ
s1ox1X0Qjzoix2y8RN0zhPLx+Iji6bZyy4a+ycu1kSIQgBp9sSTmj+0J9gJSC/0n
fAfsgcWiwutsMfkvxwTJm1DvurlK1/dOFqBDzZ6M+KGZYq1ucsBrlSu8t1iqIZ11
28FdSTMOWJ7DNCJx+FiIasILxRW65CUOnMYHiHHtpaUnm3a5Zg/SV0xnAr2OuvA/
rGj/QU6VOdtV7ti7R8QjrQJVGgtlPF5FbopbzDS9kyvBH/nigQAJCeFB6mcDbcPd
Jkiz8TzZJWo6ONPv/2+DMZXzwHglo9pXWY3RxtsJ5WayJZE2++tOvVGQTRiDlZUP
HubH0hfvy3hgdN///8Iq446Fwnof0UXVvRAqfsACbNK8zQ6ctXYP+vsNQWDlIK+r
lNpeNU+MWbewY6Qu90ezc0re6t3d76CZIyOYGETOI55Zo+C9VN5JFuz/8SAvk/th
cA+Gd6mB070MH6fOyiu/nAHzVjuMhGLV8wu+0q3sXtpoZ4TCyHZ6bboVl8di8Yxo
/cihCRL576KqOjoIwY2ZUUtVJdqWaOrsGN0mVbO7LCVoXP/F2O86QtPVOBdF+Pdo
c1siT/B6y5jw8CLB/lgKlw==
//pragma protect end_data_block
//pragma protect digest_block
0x7sEgid9tyvlIluQhBt4fqrazk=
//pragma protect end_digest_block
//pragma protect end_protected
