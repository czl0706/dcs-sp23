//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2BMfQiLIduEn12bbOTePlcXzs2ypUFChR8PV9GplvQ4BVitJOGutPNmbH39BZ8rN
trMxwrJGyhnGl8XEZ0VGnwjYPwvrhQ3UdCUNirsZahdP8Va5FQ1GZW1E+mggWE13
UVHBpm3MZPdfphp9prLT9xm5bdRH1c3/k35DtzGI2wfxyfpHHH0MXA==
//pragma protect end_key_block
//pragma protect digest_block
jM5lTFsxJIBkdhnLalEGAIrX4O8=
//pragma protect end_digest_block
//pragma protect data_block
VYtyYXx2AnNtmHKQHJ4HnsWCLmjqGSXjQRQnHiUkwdLXj+zAjuEHBt3tlIGwuQlJ
OYVRD9gNv4oljYET5KYew8O4QaG6dpoiHEKw6DMccdouALynh21omcNJ4OAq9YKs
iGHzJv+aXbYYFfEDeqiJJQ74R5Mn+6PoWKXBxL1j9JxhyntNzMFG5HRoKUh/R8m3
5fm6fLmiQdzAsYhKhAgNmXZXvpbBUIPKgDmrOlpPyhyRsLTtJiZN0lpJOmlDGujc
E60qEXuSQjr8WYD3rbTAqNs3KO3zdG4IUAsGUxGT+QvXYmP2Goho9R1YxBAhXvrn
BWTYXdp+VwcN2JjLzz5T1kMjZmhiX54PeuH1Ty+Yh9M3OfaTbFWlxVSw+Br8kFFz
IfoQxNjp7cC6KMlp7ZLh/WT5ypk7XNu28etzpc3tu1KpG/a38aOizkH81c6V/GB2
Cv8z0HiOzGHMfh4fFMI1PFO1xy+aw9Iq2Tl2b5nLv9Y9jDJDC36wxU2w1vGs6YFK
Xe3op3yhuCXO3PAThwB84NhQXmP6oDVZeaB+RhSU/7PQWKv7xo6vsTdIorwEl8V7
HBHEaAjzMbqEinUFMNgsjpQSpS0CZpBylsOuC8Un7WJoiSZ+u0wAKcp5y7XjAC7K
ONWV+IuQadV+I7Quj7+zVAAZjlECLZ/BNPRoivpvWJa+iNXvRUxk087WzTj4ZdDL
9/31rWQuksLa3RdQDs0s/ZxxIgBRr99rUaSIuNkIuG503BG65JgaB17zKpNjrGot
AQQmMQVB+yVCAty0Oc5pCRz8xdAC275foMWbID5odXNCTERyHF6/myJcgtw8Mldl
rgzAJQXNLP3aNKmINY8SzXxrEbKXdyDNJJ9JMZ6AIJpJgDx0bGOVJV0OArRehgfw
5n0uYLHFDje4QXq8eKiB6DyBN+uROHzyc4WIZfrrdHbcJ6lJSBgVjH20WG/Xt/2H
oYpKIQOXbC59++odXEsAyF0sz3rSBEhmc9yJNum/mDxkLTNppNt/BRuO/c0X40Jy
b11Fbhb5geIdTaTtD24rJaKEsXNeYTA/spkRWVCFxzX5YmTut2t2YMAn8sf4jvk5
IYtElyeONpCvjGInTE5pMWSmrawtyyuNuSCDBZqjwUDS0jZLHr22qD7yv7nF3FSf
PXYAXVK93wOH5DmpWNWHEDbKe49JiriV8fq3/u9nDmoso6ZKsUK2kQkm5oot/BkH
rKgknRSRZsgcbzE4fOcm56USKLDJk3OKUXzthNAoVHgqnjRMZpE7NAlxBK43KeLk
5gzroAhZ6LiTGY8bSIAn3qx7qpS3iAf2S+uNxkBAM0T7tRL44eWQLqCX9RvEPjlb
LGtQbJD3jwbkksTLVutnKW+n2sLIK/md0LPB+3mLJRDELGKWmR7SP5Yb+m/WYAlU
AQLs5l6GRlL13ZlFeYvajxq2xzvJn4NXKjNLtLZlXoqCAwLacfGitsVJZOyjdK6o
HGSW6L6C8g+vEcv5+fU9vIooMgeh72ysDJARTUr3EnBUpvMgjbnHStOdQsix9css
thuNdo5H2Dm0gzINgGi7jQFIbjvNpuoLyYXC2rSPz0+sDXG6cuWZYMi27fdIz1B6
+dqmchKuuKjzlEPItmzWpiyhm9xf5D0yeDD+YbuPQOCq9gaIAlpWgvzXGhFFl6ss
METD5ixB63PChc5Bcv0KqYApo22ORWn7o8fIwb/CtRS+5KzCktyd+FU8rpxSDKsK
Y2Qm9goQgta1oDWpxuCixCjQePkcvpMZvwwY47HO2LMO90eQWfFaNTHis/lkFAPF
3aAtn/aCvwsw2j9CZfDNrrG4946cfjtRtLzgUj87e820PQYhF8zJAB9My2gRJs3z
B3S/enpkhxGaLKiKkZQ8IjeUZvn4OaRi6vhuS3JFTbSfSHZFtoVkmwVm0P90pDJX
nrgsFlfpHVU9cvoiWRrmLj52KRUIXFSsiUO8TRwQaQKWoAzL85ulKjVLeaBo/gZK
gQ4X9OzxRMdEh9Sv9iDV6c83qY7a6xb1u50Wg7Vf+3K4XOdEVwQfQYHoKel+LvSp
fk3CyaFPEhNvIHt9EK5gko/cZchr8wfMQjMhhLx9XCwMY5BMxhLXM4EXws1KF2ze
c6TEmXV4hxfkOzjMAE51HfwhWFVfNpgtOMlqUpa6zfHxd5YbdXkASZxzM9DwNkOO
fLacCuicH9NDJQ22m3XZHfqMF6oBvUt11XMTXlV7rhIaILGsTlhKfuHmLAkh5Zic
eZ/VHWu7YcM3/rvU6vigly7n81t897UFrReu9S3idDR2weYsOANY2kPMBJ8xhMTN
D58Im2ZF7O390ONFi1qwfj6CxXAOISTtegJGhCoP7Eb1s1U9f0ccPB/zW37+imIg
XvsIQZOrzFI5cIJjxNIUKlNZcgcWKraRFGw37HI8fit6DRUhN7hVNjWzxOmI+Aow
gdUAm6yoVyZbDNG0GjZoM7U4VDgaMNB17Z0PzDuYq/AAUp2uPBA7SRONufmGNWhn
twTFW0FZ+xt+L3b/yFzZWQatujJsOUXsWFqO2VhnmD1dknwM4WxTPeGbxEnTMwQg
DDGhpy2UzfmtExwnK8o8ocwkjOstUb90GIK1yJCHIJE31RbSlQdBa+HRI9dRgvk4
IlmLOTASM4+II07tZVduZ6kzNoQcA0VhwKo5xKqNN98iU4qD/536pIjMSdtmV8Z0
i4BeSqOxutTxXmNinsWXIXkNqDUQIMb+7zzfnHb7g3otEB83ywTLe+n3qwKefSI2
jKysZd1m/ns3mm17r/VPBCy3P2Pix1Gjmyw52GnqgAfaCal7/NWN4rT643tbCK58
hidjRnVO9D8Wq/DVvpjyx8sn78uSu3XiY3SmYCGkHVmudoQbYfDPZWd5a3OrfY3d
rENO8at2YTXr7zxn81ACJH1r/dHVUHYBBEtwKE+vNsBLYNSulG4IZyDqzA59LwOP
zza5vS6hv5aLe0KY6s1OcTHyT/mZAj25AtHvivJMNqXUhSuVfO4gnHLuIXiePw5S
OSCxRyJ3wONlYi907kHfxsv3B7fJ+ZCDgy5bqXa1QE4Gj0RMqZkkK0jXZG5rzWva
0oQjS9yGfiE2H8y7y8+dunHSHV5lh1lDDSA3GBuk2OwYNaEte/qTFcSkM4GbG57h
Xn04nG425AfloIOrzqdwjE017Tx7qKR5SihBvQUhZreo36Czw6w1DNYDVNmyyxp4
0FEoaNFSkYXNGqk0qMcaum6AyskXUQZ6RYudUi7pa9TceHO3NHPBlYxF78PhyAoj
hr/hZiyswNRL6NVS6lWRXb1gitlrE0FRRyyrrj85+7xP7QsjHfQ4x57lHhbcRYC7
qxa9s4FycyRbsE3wjVCt1wt3J4nKDm6AxKoDrdaa36QmVsbDQw7mE2UIwLPBTz4R
GgSdjYeOlMohTj6MQ3H5YFApy93HDHY0CUF2gXD+d6ccWW5Nwt86bgPP7a/mEdM7
b1ba3GT2gJI7hfcol/+9SeMP5eas62ji3r66fK4P/sNvxOAPxMWeV8VAtzmRVMWN
ZRKaQ5tzHJA5gsGyyCn04VHKhl3pNMBEBmqGVNcdVyXPkgYtfl7xYwXWSs4qIPQY
0p0x8XvqZURD2wlE831FKDH4jJ0yXf/an9/QPWvomTj/bm9NZnOFlY3KqcRFtElh
LuhzIRBB9MgYiH9LLS+x+EquD7k/e0gCpIgy5ZLYeV9vkulFc5jGzgXiKn7n2ucx
Z9PfSU3ub7BaI3DjvYjPpEBoF5HL9De4O6F0yH1GMn9gomk/EUcfMXLE+8tyOZmI
Rj30uvkeEOXu62TvpGkaXQ4GdbkFAqwRljP0SkPjRMhX0oDF5ItgReVEUBFYEq37
oU2y+2Fk90b1vyLx2nqvQzdzlr3SCTdU3aIwN+LwXd5L58v+BY9nAWCM4eCh0zBx
ykb3m00uq3wRJ/e+uCGdZ2PWszYCliAd4qEqrY3HDPFRHhO+WEWIurnqJhIk1HiM
UCMjUR1o1KfMlWv7Buwx00me2HXhyZKyNmktvul+sSmUQ8E7EzYcJtH3VAiDFhGD
2ME6Hyhblf6P4LPwAy9hLTTCkpj2NjRdiVaxYukN8nWT2LgCMXksEvJ8cU5jytoD
Iduc2xQ2mOf4RESWcxgQP+cc2dpqWfhUATzklltl+uO5fx5hWa2Cvhic5SZuVtyi
GmU2fFTEA5vrBAjJy9WzipFM6oBanGwr5cNmft7b7wz9V9rNRlDImnkhAPhq2L37
9hITFdIBnJPYaymjjriOsjvBuq4RUeyShUZD/mJAf7D1eKc484yoUqGUlVrs2hD6
YmKFBjtHJ576mjOpEb8kkCmSS9adAa7kD2E75Qg9BxqRzOrRxKNX5z8NvW3leedP
pyHt5kymU4quvsDNkdg4iVy/v3cSlNIDu8ASwC41Jq8+oJYr0U6r28If2MBhdw03
ChA233c3SYELziqa/ZBiVAPY7V8Yn4Gq5DWaNIFZn7iswCT7+5cj/L3qlMFKkSBo
JBUZc5jRdUSX/QP8kKXVTseX2VQDpK31U/18Dz41d/vc6TodPb0LjTUKy4kgb2G3
r75M2x28U769g7Ti2CjvBzppBiXmw7+gUKFRPp8RrHoqq8wC9YtCea6RXeZnzOSw
nQT2XgC1F46VtPKSSYX4xH/gggNwUd9Z//iDRMR5c7j76PJbeorCMjxi+Enfvj8J
L089zzr3jHaa7XWkND0wPa+NcI96qwoAQRazpqDofJRo3FwReYqW6xzR33aqIvG7
qGhOJLtyteo+XniMSQZs6z6S2ZW52IZMN7vlW8Z54lDS8CzFLUtX7y4k2RrCUPtA
y6s69+kdUdkLJi9XXG68vxqE2epLeqWz/xd1w8K/tfsvTALC1EpjKsaRJ72VSlRj
6k4H6T8Z1lqifKYVBkcOXx7gima/W/pMeOetSQMTueNcR8qfaF7XdnDWdpUqa352
zo85LjYMxsweiWjvLeBOEr5lWlRHGs23qRT/KLOGAxzT8Qbc4gCExq4OXcvLg1z4
/vc8vWQCJFAUtuISMWt2hSq6dNftvFQJN5zRf/BbbTrKy1J+Ptsgvv0KTjRGjjRW
THxuqYxVxUiQ5D/DV4yXsR8V5ApOjw0fDFTR3E5E++5TKQcqeiMIRffG78jSiquS
sgcS5bvWn1PWRNKMsKje7BzdWayQ36OjpRPEzXgNIldEqbKu3mHJiQgSaZ5YVOGi
Ij2qirhQPAVK5Znu8yo11+7BWd0oyfoEjhQ+ZMfhigXalL9LkOVQ4+vui7c7Jl3X
jDz9E2vDv7W1rzgeZzfXuvVPTqDUFSrVZ0VxdUs+fUfahm+4CcDpnctbGFqNYWZy
PO0EmFspm0XbRba78c3/crF8A7SLOYIIwavIpAaAaypYtZZBesduzdO3m3Wfe8T6
IDKtDCeYvALG5qVKob/JONiaXPQCtQnXy9deQ3w9I4XWMFbTvufcd1NeryFyUOGQ
3DpgmYFoyPTGcFTGUejbKsM2z2rj6iQJ0wC4g9zMwmkvJdg/aK+wndOQiXRwDFgU
Zw9hlzyoUjAkxUYBcmW0UefhEQ5+/BR5g/byFNxU4B4kLxS2s/aQcEfNHNwh4vxm
ZaPfC6zPt9vyn4SK8JaVfj3WJhuF6h6nuMldqmSg5BmgH48gMgQQek0hcOX29/Fs
c9Tyhu0Yxyk4ESHbMATZYuT+/zbC3ka9D9P3YFL/BGYd0dpAjyS6J7Eg9SwyA+36
snswv1sh5S1CApnEQIiIkWtsVNhglbVNkSDCWPBgADQKq/wSGnUONkISMgPOaDEO
SP12Re6OwRfOaVRUMpaSzCWJ6po5afoXLir3o4EiOcuqKfXKV9odpz8KYYdak4rF
G3uOlOshe6fSFUJZnqOPSkMgefUT9+Jk9GKt7ZW2gbEQvTwbpREJ/l7U6g36hYBI
sGxL6EOn8QpqBT4pSOcznnhdhQ8PR8b/GddPtKaNZOExRHRwDqJ6uRkunhgstE40
0voIxCNoJROvU4OPZQx8lPK81gJxoYeT7Eq7OAZm7/3SpWbXovpmCPSiktzpuY7c
jR52X2b81InZz4PtYqrrjp6zIWk8Psgb8tIl3cwwXWYbVy1OdoN4fbVFyrQG3C7b
WG9FMr6VpKIYqf4RV/ZvC6amA2JHh5xMVTud1xNm1D4xEOkYEkf4QAGEEkrFmETG
sO4XvW2BOMLo/bqal883Heq1705Rt2Mri4NiLwjNKihAV865TvX9KzuwQTOOQUlA
hmZZu7cQZBuIcpiE3dS49g4NGa7ph/M2rgJMOJhMQ6ENLmVtAHi90D7Ab/L/A+Rp
xhfIrquolvxZP7IwKwlrx3ZlO9FUXqbWVqzWSD96jz9qrtXm/N5dGQ2eMTgbuRcl
gSRAziIrb1d72SnJlvg21Mu5o4xKS5Z9dZzeB+7V1ZHAH6WAu4VdtPnT7/RWy98R
btKSHv5iSwYFWFT2PwuiZpp3ymoa0bxyvtayAntq0iaLXnJnZEcAbFY9afLslZWm
lBEJDg6nEortPwYY208sNvI6cqob6VXhHUk9CgsnilnndPpKQ5EUhHzOw/9j8f9z
lnR2OhqDtwzw4L1u7wEvKLa2Nqjx50MtaHzJdNxsAF4LDmuZDKhyiiQOcXBFlUpU
rYzzx8Qlo8aTRM8GKllUOR1sXJvZ74m+0k7HxtW/yVSTHFsy27aewl95LDFngqzo
HhRB4Ia9IoMw/uQanaVAKewcS87CuOpvLpNH9th7msj5GHeG1sHHzvEIizpWmRS0
Q772PtmuUdux9DneYkEaCOGozsOBSI7IvTPhtmBYJqn0AjPDOnvCQmvlNJLElwea
+1TTydQ4Aw1mAMaIRNeZq6nqXrHnnfh+khm6kZFZ4Y+kELMx3cBB6lzwpA9UBZ9D
E2x6yFX1wRjFZtZWpDrbGv0i23JQi66lFQj7VM+033w9p7HmQCGV7493A/U4yM5s
BPNUf3sENDRNhcDOCUdLEDCJ+ofX+3pIrza/3umHNx/u4lgQ0z0zjzCcYevs7i+6
VousBhNruZFUO4IQ39BFqbjbJQZaEu0DO0EPdkOXDFUXDh/JogEWBEmXWA+9p0jr
rajaXxq2diRKSGVGGCySHd4h0/ybRUu4xsL4A4KVHacDuWQblBFJJoh9RSb32rCb
P59iPxSZepA/HqoItEkXhoiHo87HRUOGsb3aOekoTLkU1Js6SBYK3OY30rVp2dPZ
wP3vsrq8vt3aIX3WIcSmHJfSO7Iq3mn/VbHmGcZ7UtCVrC8JFcV8RK/nDcWeFoV0
iKQDYefC3orWHALrfnVhMgc20W+Nn6qFxlTQrfdocSQ=
//pragma protect end_data_block
//pragma protect digest_block
5D/h+wNGg9SgjpObVWXUfHnUrMM=
//pragma protect end_digest_block
//pragma protect end_protected
